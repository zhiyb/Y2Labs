// D1 - model solution
// registers C and AQ, code as suggested in the briefing lecture
/*
   author: tjk
   last revision: 17 Oct' 13
*/

module register #(parameter n = 4)
				(input logic clock, reset, add_shift, shift, C,
				 input logic[n - 1:0] Qin, Sum, output logic[n * 2 - 1:0] AQ);

logic Creg; // MSB carry bit storage

always_ff @ (posedge clock)
  if (reset)  // clear C,A and load Q
  begin
   Creg <= 0;
   AQ[n * 2 - 1:n] <= 0;
   AQ[n - 1:0] <= Qin; // load multiplier into Q
  end
  else if (add_shift) // add, then shift
   {Creg,AQ} <= {1'b0,C,Sum,AQ[n - 1:1]};
  else if (shift) // shift A, Q
   {Creg,AQ} <= {1'b0,Creg,AQ[n * 2 - 1:1]};
endmodule
