// Verilog test bench for D2 chip design

`timescale 1ns/1ps

module test_TEAMJ_Adder_DESIGN;

// declare DUT input signals as "reg"
// declare DUT output signals as "wire"

reg A3;
reg A4;
reg A5;
reg A6;
reg A7;
reg A8;
reg A9;
reg A10;
reg A11;
wire Q3;
wire Q4;
wire Q5;
wire Q6;
wire Q7;
integer errors_Q3;
integer errors_Q4;
integer errors_Q5;
integer errors_Q6;
integer errors_Q7;

// declare error count

integer errors;

// instance Device Under Test
//   assumes top-level OrCAD schematic is named "TEAMJ_Adder_DESIGN"

`ifdef DUT
  `DUT DUT(
`else
  TEAMJ_DESIGN DUT(
`endif
   .A3(A3),
   .A4(A4),
   .A5(A5),
   .A6(A6),
   .A7(A7),
   .A8(A8),
   .A9(A9),
   .A10(A10),
   .A11(A11),
   .Q3(Q3),
   .Q4(Q4),
   .Q5(Q5),
   .Q6(Q6),
   .Q7(Q7)
);

// monitor the I/O
initial
  begin
    $display( "Simulation Begins" );
    $display ( "  AAAAAAAAA  QQQQQ" );
    $display ( "  345678911  34567" );
    $display ( "         01       " );
    $display ( "                  " );
    `ifdef no_monitor
    `else
    $monitor ( "  ",
      A3,
      A4,
      A5,
      A6,
      A7,
      A8,
      A9,
      A10,
      A11,
      "  ",
      Q3,
      Q4,
      Q5,
      Q6,
      Q7,
      "  @ %d ns", $time   );
    `endif
  end

// stimulii

initial
  begin
    errors = 0;
    errors_Q3 = 0;
    errors_Q4 = 0;
    errors_Q5 = 0;
    errors_Q6 = 0;
    errors_Q7 = 0;
    $display ( "v 000000000  00000");
    apply_vector ( 9'b000000000,5'b00000,
                   9'b111111111,5'b11111);
    $display ( "v 000001000  10000");
    apply_vector ( 9'b000001000,5'b10000,
                   9'b111111111,5'b11111);
    $display ( "v 000000100  01000");
    apply_vector ( 9'b000000100,5'b01000,
                   9'b111111111,5'b11111);
    $display ( "v 000001100  11000");
    apply_vector ( 9'b000001100,5'b11000,
                   9'b111111111,5'b11111);
    $display ( "v 000000010  00100");
    apply_vector ( 9'b000000010,5'b00100,
                   9'b111111111,5'b11111);
    $display ( "v 000001010  10100");
    apply_vector ( 9'b000001010,5'b10100,
                   9'b111111111,5'b11111);
    $display ( "v 000000110  01100");
    apply_vector ( 9'b000000110,5'b01100,
                   9'b111111111,5'b11111);
    $display ( "v 000001110  11100");
    apply_vector ( 9'b000001110,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 000000001  00010");
    apply_vector ( 9'b000000001,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 000001001  10010");
    apply_vector ( 9'b000001001,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 000000101  01010");
    apply_vector ( 9'b000000101,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 000001101  11010");
    apply_vector ( 9'b000001101,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 000000011  00110");
    apply_vector ( 9'b000000011,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 000001011  10110");
    apply_vector ( 9'b000001011,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 000000111  01110");
    apply_vector ( 9'b000000111,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 000001111  11110");
    apply_vector ( 9'b000001111,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 010000000  10000");
    apply_vector ( 9'b010000000,5'b10000,
                   9'b111111111,5'b11111);
    $display ( "v 010001000  01000");
    apply_vector ( 9'b010001000,5'b01000,
                   9'b111111111,5'b11111);
    $display ( "v 010000100  11000");
    apply_vector ( 9'b010000100,5'b11000,
                   9'b111111111,5'b11111);
    $display ( "v 010001100  00100");
    apply_vector ( 9'b010001100,5'b00100,
                   9'b111111111,5'b11111);
    $display ( "v 010000010  10100");
    apply_vector ( 9'b010000010,5'b10100,
                   9'b111111111,5'b11111);
    $display ( "v 010001010  01100");
    apply_vector ( 9'b010001010,5'b01100,
                   9'b111111111,5'b11111);
    $display ( "v 010000110  11100");
    apply_vector ( 9'b010000110,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 010001110  00010");
    apply_vector ( 9'b010001110,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 010000001  10010");
    apply_vector ( 9'b010000001,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 010001001  01010");
    apply_vector ( 9'b010001001,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 010000101  11010");
    apply_vector ( 9'b010000101,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 010001101  00110");
    apply_vector ( 9'b010001101,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 010000011  10110");
    apply_vector ( 9'b010000011,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 010001011  01110");
    apply_vector ( 9'b010001011,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 010000111  11110");
    apply_vector ( 9'b010000111,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 010001111  00001");
    apply_vector ( 9'b010001111,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 001000000  01000");
    apply_vector ( 9'b001000000,5'b01000,
                   9'b111111111,5'b11111);
    $display ( "v 001001000  11000");
    apply_vector ( 9'b001001000,5'b11000,
                   9'b111111111,5'b11111);
    $display ( "v 001000100  00100");
    apply_vector ( 9'b001000100,5'b00100,
                   9'b111111111,5'b11111);
    $display ( "v 001001100  10100");
    apply_vector ( 9'b001001100,5'b10100,
                   9'b111111111,5'b11111);
    $display ( "v 001000010  01100");
    apply_vector ( 9'b001000010,5'b01100,
                   9'b111111111,5'b11111);
    $display ( "v 001001010  11100");
    apply_vector ( 9'b001001010,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 001000110  00010");
    apply_vector ( 9'b001000110,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 001001110  10010");
    apply_vector ( 9'b001001110,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 001000001  01010");
    apply_vector ( 9'b001000001,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 001001001  11010");
    apply_vector ( 9'b001001001,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 001000101  00110");
    apply_vector ( 9'b001000101,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 001001101  10110");
    apply_vector ( 9'b001001101,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 001000011  01110");
    apply_vector ( 9'b001000011,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 001001011  11110");
    apply_vector ( 9'b001001011,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 001000111  00001");
    apply_vector ( 9'b001000111,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 001001111  10001");
    apply_vector ( 9'b001001111,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 011000000  11000");
    apply_vector ( 9'b011000000,5'b11000,
                   9'b111111111,5'b11111);
    $display ( "v 011001000  00100");
    apply_vector ( 9'b011001000,5'b00100,
                   9'b111111111,5'b11111);
    $display ( "v 011000100  10100");
    apply_vector ( 9'b011000100,5'b10100,
                   9'b111111111,5'b11111);
    $display ( "v 011001100  01100");
    apply_vector ( 9'b011001100,5'b01100,
                   9'b111111111,5'b11111);
    $display ( "v 011000010  11100");
    apply_vector ( 9'b011000010,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 011001010  00010");
    apply_vector ( 9'b011001010,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 011000110  10010");
    apply_vector ( 9'b011000110,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 011001110  01010");
    apply_vector ( 9'b011001110,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 011000001  11010");
    apply_vector ( 9'b011000001,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 011001001  00110");
    apply_vector ( 9'b011001001,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 011000101  10110");
    apply_vector ( 9'b011000101,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 011001101  01110");
    apply_vector ( 9'b011001101,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 011000011  11110");
    apply_vector ( 9'b011000011,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 011001011  00001");
    apply_vector ( 9'b011001011,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 011000111  10001");
    apply_vector ( 9'b011000111,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 011001111  01001");
    apply_vector ( 9'b011001111,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 000100000  00100");
    apply_vector ( 9'b000100000,5'b00100,
                   9'b111111111,5'b11111);
    $display ( "v 000101000  10100");
    apply_vector ( 9'b000101000,5'b10100,
                   9'b111111111,5'b11111);
    $display ( "v 000100100  01100");
    apply_vector ( 9'b000100100,5'b01100,
                   9'b111111111,5'b11111);
    $display ( "v 000101100  11100");
    apply_vector ( 9'b000101100,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 000100010  00010");
    apply_vector ( 9'b000100010,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 000101010  10010");
    apply_vector ( 9'b000101010,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 000100110  01010");
    apply_vector ( 9'b000100110,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 000101110  11010");
    apply_vector ( 9'b000101110,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 000100001  00110");
    apply_vector ( 9'b000100001,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 000101001  10110");
    apply_vector ( 9'b000101001,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 000100101  01110");
    apply_vector ( 9'b000100101,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 000101101  11110");
    apply_vector ( 9'b000101101,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 000100011  00001");
    apply_vector ( 9'b000100011,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 000101011  10001");
    apply_vector ( 9'b000101011,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 000100111  01001");
    apply_vector ( 9'b000100111,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 000101111  11001");
    apply_vector ( 9'b000101111,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 010100000  10100");
    apply_vector ( 9'b010100000,5'b10100,
                   9'b111111111,5'b11111);
    $display ( "v 010101000  01100");
    apply_vector ( 9'b010101000,5'b01100,
                   9'b111111111,5'b11111);
    $display ( "v 010100100  11100");
    apply_vector ( 9'b010100100,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 010101100  00010");
    apply_vector ( 9'b010101100,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 010100010  10010");
    apply_vector ( 9'b010100010,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 010101010  01010");
    apply_vector ( 9'b010101010,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 010100110  11010");
    apply_vector ( 9'b010100110,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 010101110  00110");
    apply_vector ( 9'b010101110,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 010100001  10110");
    apply_vector ( 9'b010100001,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 010101001  01110");
    apply_vector ( 9'b010101001,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 010100101  11110");
    apply_vector ( 9'b010100101,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 010101101  00001");
    apply_vector ( 9'b010101101,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 010100011  10001");
    apply_vector ( 9'b010100011,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 010101011  01001");
    apply_vector ( 9'b010101011,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 010100111  11001");
    apply_vector ( 9'b010100111,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 010101111  00101");
    apply_vector ( 9'b010101111,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 001100000  01100");
    apply_vector ( 9'b001100000,5'b01100,
                   9'b111111111,5'b11111);
    $display ( "v 001101000  11100");
    apply_vector ( 9'b001101000,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 001100100  00010");
    apply_vector ( 9'b001100100,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 001101100  10010");
    apply_vector ( 9'b001101100,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 001100010  01010");
    apply_vector ( 9'b001100010,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 001101010  11010");
    apply_vector ( 9'b001101010,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 001100110  00110");
    apply_vector ( 9'b001100110,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 001101110  10110");
    apply_vector ( 9'b001101110,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 001100001  01110");
    apply_vector ( 9'b001100001,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 001101001  11110");
    apply_vector ( 9'b001101001,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 001100101  00001");
    apply_vector ( 9'b001100101,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 001101101  10001");
    apply_vector ( 9'b001101101,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 001100011  01001");
    apply_vector ( 9'b001100011,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 001101011  11001");
    apply_vector ( 9'b001101011,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 001100111  00101");
    apply_vector ( 9'b001100111,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 001101111  10101");
    apply_vector ( 9'b001101111,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 011100000  11100");
    apply_vector ( 9'b011100000,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 011101000  00010");
    apply_vector ( 9'b011101000,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 011100100  10010");
    apply_vector ( 9'b011100100,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 011101100  01010");
    apply_vector ( 9'b011101100,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 011100010  11010");
    apply_vector ( 9'b011100010,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 011101010  00110");
    apply_vector ( 9'b011101010,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 011100110  10110");
    apply_vector ( 9'b011100110,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 011101110  01110");
    apply_vector ( 9'b011101110,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 011100001  11110");
    apply_vector ( 9'b011100001,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 011101001  00001");
    apply_vector ( 9'b011101001,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 011100101  10001");
    apply_vector ( 9'b011100101,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 011101101  01001");
    apply_vector ( 9'b011101101,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 011100011  11001");
    apply_vector ( 9'b011100011,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 011101011  00101");
    apply_vector ( 9'b011101011,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 011100111  10101");
    apply_vector ( 9'b011100111,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 011101111  01101");
    apply_vector ( 9'b011101111,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 000010000  00010");
    apply_vector ( 9'b000010000,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 000011000  10010");
    apply_vector ( 9'b000011000,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 000010100  01010");
    apply_vector ( 9'b000010100,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 000011100  11010");
    apply_vector ( 9'b000011100,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 000010010  00110");
    apply_vector ( 9'b000010010,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 000011010  10110");
    apply_vector ( 9'b000011010,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 000010110  01110");
    apply_vector ( 9'b000010110,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 000011110  11110");
    apply_vector ( 9'b000011110,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 000010001  00001");
    apply_vector ( 9'b000010001,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 000011001  10001");
    apply_vector ( 9'b000011001,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 000010101  01001");
    apply_vector ( 9'b000010101,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 000011101  11001");
    apply_vector ( 9'b000011101,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 000010011  00101");
    apply_vector ( 9'b000010011,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 000011011  10101");
    apply_vector ( 9'b000011011,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 000010111  01101");
    apply_vector ( 9'b000010111,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 000011111  11101");
    apply_vector ( 9'b000011111,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 010010000  10010");
    apply_vector ( 9'b010010000,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 010011000  01010");
    apply_vector ( 9'b010011000,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 010010100  11010");
    apply_vector ( 9'b010010100,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 010011100  00110");
    apply_vector ( 9'b010011100,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 010010010  10110");
    apply_vector ( 9'b010010010,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 010011010  01110");
    apply_vector ( 9'b010011010,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 010010110  11110");
    apply_vector ( 9'b010010110,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 010011110  00001");
    apply_vector ( 9'b010011110,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 010010001  10001");
    apply_vector ( 9'b010010001,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 010011001  01001");
    apply_vector ( 9'b010011001,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 010010101  11001");
    apply_vector ( 9'b010010101,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 010011101  00101");
    apply_vector ( 9'b010011101,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 010010011  10101");
    apply_vector ( 9'b010010011,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 010011011  01101");
    apply_vector ( 9'b010011011,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 010010111  11101");
    apply_vector ( 9'b010010111,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 010011111  00011");
    apply_vector ( 9'b010011111,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 001010000  01010");
    apply_vector ( 9'b001010000,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 001011000  11010");
    apply_vector ( 9'b001011000,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 001010100  00110");
    apply_vector ( 9'b001010100,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 001011100  10110");
    apply_vector ( 9'b001011100,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 001010010  01110");
    apply_vector ( 9'b001010010,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 001011010  11110");
    apply_vector ( 9'b001011010,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 001010110  00001");
    apply_vector ( 9'b001010110,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 001011110  10001");
    apply_vector ( 9'b001011110,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 001010001  01001");
    apply_vector ( 9'b001010001,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 001011001  11001");
    apply_vector ( 9'b001011001,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 001010101  00101");
    apply_vector ( 9'b001010101,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 001011101  10101");
    apply_vector ( 9'b001011101,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 001010011  01101");
    apply_vector ( 9'b001010011,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 001011011  11101");
    apply_vector ( 9'b001011011,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 001010111  00011");
    apply_vector ( 9'b001010111,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 001011111  10011");
    apply_vector ( 9'b001011111,5'b10011,
                   9'b111111111,5'b11111);
    $display ( "v 011010000  11010");
    apply_vector ( 9'b011010000,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 011011000  00110");
    apply_vector ( 9'b011011000,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 011010100  10110");
    apply_vector ( 9'b011010100,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 011011100  01110");
    apply_vector ( 9'b011011100,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 011010010  11110");
    apply_vector ( 9'b011010010,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 011011010  00001");
    apply_vector ( 9'b011011010,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 011010110  10001");
    apply_vector ( 9'b011010110,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 011011110  01001");
    apply_vector ( 9'b011011110,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 011010001  11001");
    apply_vector ( 9'b011010001,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 011011001  00101");
    apply_vector ( 9'b011011001,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 011010101  10101");
    apply_vector ( 9'b011010101,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 011011101  01101");
    apply_vector ( 9'b011011101,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 011010011  11101");
    apply_vector ( 9'b011010011,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 011011011  00011");
    apply_vector ( 9'b011011011,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 011010111  10011");
    apply_vector ( 9'b011010111,5'b10011,
                   9'b111111111,5'b11111);
    $display ( "v 011011111  01011");
    apply_vector ( 9'b011011111,5'b01011,
                   9'b111111111,5'b11111);
    $display ( "v 000110000  00110");
    apply_vector ( 9'b000110000,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 000111000  10110");
    apply_vector ( 9'b000111000,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 000110100  01110");
    apply_vector ( 9'b000110100,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 000111100  11110");
    apply_vector ( 9'b000111100,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 000110010  00001");
    apply_vector ( 9'b000110010,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 000111010  10001");
    apply_vector ( 9'b000111010,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 000110110  01001");
    apply_vector ( 9'b000110110,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 000111110  11001");
    apply_vector ( 9'b000111110,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 000110001  00101");
    apply_vector ( 9'b000110001,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 000111001  10101");
    apply_vector ( 9'b000111001,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 000110101  01101");
    apply_vector ( 9'b000110101,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 000111101  11101");
    apply_vector ( 9'b000111101,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 000110011  00011");
    apply_vector ( 9'b000110011,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 000111011  10011");
    apply_vector ( 9'b000111011,5'b10011,
                   9'b111111111,5'b11111);
    $display ( "v 000110111  01011");
    apply_vector ( 9'b000110111,5'b01011,
                   9'b111111111,5'b11111);
    $display ( "v 000111111  11011");
    apply_vector ( 9'b000111111,5'b11011,
                   9'b111111111,5'b11111);
    $display ( "v 010110000  10110");
    apply_vector ( 9'b010110000,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 010111000  01110");
    apply_vector ( 9'b010111000,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 010110100  11110");
    apply_vector ( 9'b010110100,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 010111100  00001");
    apply_vector ( 9'b010111100,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 010110010  10001");
    apply_vector ( 9'b010110010,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 010111010  01001");
    apply_vector ( 9'b010111010,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 010110110  11001");
    apply_vector ( 9'b010110110,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 010111110  00101");
    apply_vector ( 9'b010111110,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 010110001  10101");
    apply_vector ( 9'b010110001,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 010111001  01101");
    apply_vector ( 9'b010111001,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 010110101  11101");
    apply_vector ( 9'b010110101,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 010111101  00011");
    apply_vector ( 9'b010111101,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 010110011  10011");
    apply_vector ( 9'b010110011,5'b10011,
                   9'b111111111,5'b11111);
    $display ( "v 010111011  01011");
    apply_vector ( 9'b010111011,5'b01011,
                   9'b111111111,5'b11111);
    $display ( "v 010110111  11011");
    apply_vector ( 9'b010110111,5'b11011,
                   9'b111111111,5'b11111);
    $display ( "v 010111111  00111");
    apply_vector ( 9'b010111111,5'b00111,
                   9'b111111111,5'b11111);
    $display ( "v 001110000  01110");
    apply_vector ( 9'b001110000,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 001111000  11110");
    apply_vector ( 9'b001111000,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 001110100  00001");
    apply_vector ( 9'b001110100,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 001111100  10001");
    apply_vector ( 9'b001111100,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 001110010  01001");
    apply_vector ( 9'b001110010,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 001111010  11001");
    apply_vector ( 9'b001111010,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 001110110  00101");
    apply_vector ( 9'b001110110,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 001111110  10101");
    apply_vector ( 9'b001111110,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 001110001  01101");
    apply_vector ( 9'b001110001,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 001111001  11101");
    apply_vector ( 9'b001111001,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 001110101  00011");
    apply_vector ( 9'b001110101,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 001111101  10011");
    apply_vector ( 9'b001111101,5'b10011,
                   9'b111111111,5'b11111);
    $display ( "v 001110011  01011");
    apply_vector ( 9'b001110011,5'b01011,
                   9'b111111111,5'b11111);
    $display ( "v 001111011  11011");
    apply_vector ( 9'b001111011,5'b11011,
                   9'b111111111,5'b11111);
    $display ( "v 001110111  00111");
    apply_vector ( 9'b001110111,5'b00111,
                   9'b111111111,5'b11111);
    $display ( "v 001111111  10111");
    apply_vector ( 9'b001111111,5'b10111,
                   9'b111111111,5'b11111);
    $display ( "v 011110000  11110");
    apply_vector ( 9'b011110000,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 011111000  00001");
    apply_vector ( 9'b011111000,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 011110100  10001");
    apply_vector ( 9'b011110100,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 011111100  01001");
    apply_vector ( 9'b011111100,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 011110010  11001");
    apply_vector ( 9'b011110010,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 011111010  00101");
    apply_vector ( 9'b011111010,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 011110110  10101");
    apply_vector ( 9'b011110110,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 011111110  01101");
    apply_vector ( 9'b011111110,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 011110001  11101");
    apply_vector ( 9'b011110001,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 011111001  00011");
    apply_vector ( 9'b011111001,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 011110101  10011");
    apply_vector ( 9'b011110101,5'b10011,
                   9'b111111111,5'b11111);
    $display ( "v 011111101  01011");
    apply_vector ( 9'b011111101,5'b01011,
                   9'b111111111,5'b11111);
    $display ( "v 011110011  11011");
    apply_vector ( 9'b011110011,5'b11011,
                   9'b111111111,5'b11111);
    $display ( "v 011111011  00111");
    apply_vector ( 9'b011111011,5'b00111,
                   9'b111111111,5'b11111);
    $display ( "v 011110111  10111");
    apply_vector ( 9'b011110111,5'b10111,
                   9'b111111111,5'b11111);
    $display ( "v 011111111  01111");
    apply_vector ( 9'b011111111,5'b01111,
                   9'b111111111,5'b11111);
    $display ( "v 100000000  10000");
    apply_vector ( 9'b100000000,5'b10000,
                   9'b111111111,5'b11111);
    $display ( "v 100001000  01000");
    apply_vector ( 9'b100001000,5'b01000,
                   9'b111111111,5'b11111);
    $display ( "v 100000100  11000");
    apply_vector ( 9'b100000100,5'b11000,
                   9'b111111111,5'b11111);
    $display ( "v 100001100  00100");
    apply_vector ( 9'b100001100,5'b00100,
                   9'b111111111,5'b11111);
    $display ( "v 100000010  10100");
    apply_vector ( 9'b100000010,5'b10100,
                   9'b111111111,5'b11111);
    $display ( "v 100001010  01100");
    apply_vector ( 9'b100001010,5'b01100,
                   9'b111111111,5'b11111);
    $display ( "v 100000110  11100");
    apply_vector ( 9'b100000110,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 100001110  00010");
    apply_vector ( 9'b100001110,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 100000001  10010");
    apply_vector ( 9'b100000001,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 100001001  01010");
    apply_vector ( 9'b100001001,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 100000101  11010");
    apply_vector ( 9'b100000101,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 100001101  00110");
    apply_vector ( 9'b100001101,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 100000011  10110");
    apply_vector ( 9'b100000011,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 100001011  01110");
    apply_vector ( 9'b100001011,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 100000111  11110");
    apply_vector ( 9'b100000111,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 100001111  00001");
    apply_vector ( 9'b100001111,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 110000000  01000");
    apply_vector ( 9'b110000000,5'b01000,
                   9'b111111111,5'b11111);
    $display ( "v 110001000  11000");
    apply_vector ( 9'b110001000,5'b11000,
                   9'b111111111,5'b11111);
    $display ( "v 110000100  00100");
    apply_vector ( 9'b110000100,5'b00100,
                   9'b111111111,5'b11111);
    $display ( "v 110001100  10100");
    apply_vector ( 9'b110001100,5'b10100,
                   9'b111111111,5'b11111);
    $display ( "v 110000010  01100");
    apply_vector ( 9'b110000010,5'b01100,
                   9'b111111111,5'b11111);
    $display ( "v 110001010  11100");
    apply_vector ( 9'b110001010,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 110000110  00010");
    apply_vector ( 9'b110000110,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 110001110  10010");
    apply_vector ( 9'b110001110,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 110000001  01010");
    apply_vector ( 9'b110000001,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 110001001  11010");
    apply_vector ( 9'b110001001,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 110000101  00110");
    apply_vector ( 9'b110000101,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 110001101  10110");
    apply_vector ( 9'b110001101,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 110000011  01110");
    apply_vector ( 9'b110000011,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 110001011  11110");
    apply_vector ( 9'b110001011,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 110000111  00001");
    apply_vector ( 9'b110000111,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 110001111  10001");
    apply_vector ( 9'b110001111,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 101000000  11000");
    apply_vector ( 9'b101000000,5'b11000,
                   9'b111111111,5'b11111);
    $display ( "v 101001000  00100");
    apply_vector ( 9'b101001000,5'b00100,
                   9'b111111111,5'b11111);
    $display ( "v 101000100  10100");
    apply_vector ( 9'b101000100,5'b10100,
                   9'b111111111,5'b11111);
    $display ( "v 101001100  01100");
    apply_vector ( 9'b101001100,5'b01100,
                   9'b111111111,5'b11111);
    $display ( "v 101000010  11100");
    apply_vector ( 9'b101000010,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 101001010  00010");
    apply_vector ( 9'b101001010,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 101000110  10010");
    apply_vector ( 9'b101000110,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 101001110  01010");
    apply_vector ( 9'b101001110,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 101000001  11010");
    apply_vector ( 9'b101000001,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 101001001  00110");
    apply_vector ( 9'b101001001,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 101000101  10110");
    apply_vector ( 9'b101000101,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 101001101  01110");
    apply_vector ( 9'b101001101,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 101000011  11110");
    apply_vector ( 9'b101000011,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 101001011  00001");
    apply_vector ( 9'b101001011,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 101000111  10001");
    apply_vector ( 9'b101000111,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 101001111  01001");
    apply_vector ( 9'b101001111,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 111000000  00100");
    apply_vector ( 9'b111000000,5'b00100,
                   9'b111111111,5'b11111);
    $display ( "v 111001000  10100");
    apply_vector ( 9'b111001000,5'b10100,
                   9'b111111111,5'b11111);
    $display ( "v 111000100  01100");
    apply_vector ( 9'b111000100,5'b01100,
                   9'b111111111,5'b11111);
    $display ( "v 111001100  11100");
    apply_vector ( 9'b111001100,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 111000010  00010");
    apply_vector ( 9'b111000010,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 111001010  10010");
    apply_vector ( 9'b111001010,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 111000110  01010");
    apply_vector ( 9'b111000110,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 111001110  11010");
    apply_vector ( 9'b111001110,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 111000001  00110");
    apply_vector ( 9'b111000001,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 111001001  10110");
    apply_vector ( 9'b111001001,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 111000101  01110");
    apply_vector ( 9'b111000101,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 111001101  11110");
    apply_vector ( 9'b111001101,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 111000011  00001");
    apply_vector ( 9'b111000011,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 111001011  10001");
    apply_vector ( 9'b111001011,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 111000111  01001");
    apply_vector ( 9'b111000111,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 111001111  11001");
    apply_vector ( 9'b111001111,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 100100000  10100");
    apply_vector ( 9'b100100000,5'b10100,
                   9'b111111111,5'b11111);
    $display ( "v 100101000  01100");
    apply_vector ( 9'b100101000,5'b01100,
                   9'b111111111,5'b11111);
    $display ( "v 100100100  11100");
    apply_vector ( 9'b100100100,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 100101100  00010");
    apply_vector ( 9'b100101100,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 100100010  10010");
    apply_vector ( 9'b100100010,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 100101010  01010");
    apply_vector ( 9'b100101010,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 100100110  11010");
    apply_vector ( 9'b100100110,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 100101110  00110");
    apply_vector ( 9'b100101110,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 100100001  10110");
    apply_vector ( 9'b100100001,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 100101001  01110");
    apply_vector ( 9'b100101001,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 100100101  11110");
    apply_vector ( 9'b100100101,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 100101101  00001");
    apply_vector ( 9'b100101101,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 100100011  10001");
    apply_vector ( 9'b100100011,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 100101011  01001");
    apply_vector ( 9'b100101011,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 100100111  11001");
    apply_vector ( 9'b100100111,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 100101111  00101");
    apply_vector ( 9'b100101111,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 110100000  01100");
    apply_vector ( 9'b110100000,5'b01100,
                   9'b111111111,5'b11111);
    $display ( "v 110101000  11100");
    apply_vector ( 9'b110101000,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 110100100  00010");
    apply_vector ( 9'b110100100,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 110101100  10010");
    apply_vector ( 9'b110101100,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 110100010  01010");
    apply_vector ( 9'b110100010,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 110101010  11010");
    apply_vector ( 9'b110101010,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 110100110  00110");
    apply_vector ( 9'b110100110,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 110101110  10110");
    apply_vector ( 9'b110101110,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 110100001  01110");
    apply_vector ( 9'b110100001,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 110101001  11110");
    apply_vector ( 9'b110101001,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 110100101  00001");
    apply_vector ( 9'b110100101,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 110101101  10001");
    apply_vector ( 9'b110101101,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 110100011  01001");
    apply_vector ( 9'b110100011,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 110101011  11001");
    apply_vector ( 9'b110101011,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 110100111  00101");
    apply_vector ( 9'b110100111,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 110101111  10101");
    apply_vector ( 9'b110101111,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 101100000  11100");
    apply_vector ( 9'b101100000,5'b11100,
                   9'b111111111,5'b11111);
    $display ( "v 101101000  00010");
    apply_vector ( 9'b101101000,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 101100100  10010");
    apply_vector ( 9'b101100100,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 101101100  01010");
    apply_vector ( 9'b101101100,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 101100010  11010");
    apply_vector ( 9'b101100010,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 101101010  00110");
    apply_vector ( 9'b101101010,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 101100110  10110");
    apply_vector ( 9'b101100110,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 101101110  01110");
    apply_vector ( 9'b101101110,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 101100001  11110");
    apply_vector ( 9'b101100001,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 101101001  00001");
    apply_vector ( 9'b101101001,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 101100101  10001");
    apply_vector ( 9'b101100101,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 101101101  01001");
    apply_vector ( 9'b101101101,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 101100011  11001");
    apply_vector ( 9'b101100011,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 101101011  00101");
    apply_vector ( 9'b101101011,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 101100111  10101");
    apply_vector ( 9'b101100111,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 101101111  01101");
    apply_vector ( 9'b101101111,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 111100000  00010");
    apply_vector ( 9'b111100000,5'b00010,
                   9'b111111111,5'b11111);
    $display ( "v 111101000  10010");
    apply_vector ( 9'b111101000,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 111100100  01010");
    apply_vector ( 9'b111100100,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 111101100  11010");
    apply_vector ( 9'b111101100,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 111100010  00110");
    apply_vector ( 9'b111100010,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 111101010  10110");
    apply_vector ( 9'b111101010,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 111100110  01110");
    apply_vector ( 9'b111100110,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 111101110  11110");
    apply_vector ( 9'b111101110,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 111100001  00001");
    apply_vector ( 9'b111100001,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 111101001  10001");
    apply_vector ( 9'b111101001,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 111100101  01001");
    apply_vector ( 9'b111100101,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 111101101  11001");
    apply_vector ( 9'b111101101,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 111100011  00101");
    apply_vector ( 9'b111100011,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 111101011  10101");
    apply_vector ( 9'b111101011,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 111100111  01101");
    apply_vector ( 9'b111100111,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 111101111  11101");
    apply_vector ( 9'b111101111,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 100010000  10010");
    apply_vector ( 9'b100010000,5'b10010,
                   9'b111111111,5'b11111);
    $display ( "v 100011000  01010");
    apply_vector ( 9'b100011000,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 100010100  11010");
    apply_vector ( 9'b100010100,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 100011100  00110");
    apply_vector ( 9'b100011100,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 100010010  10110");
    apply_vector ( 9'b100010010,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 100011010  01110");
    apply_vector ( 9'b100011010,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 100010110  11110");
    apply_vector ( 9'b100010110,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 100011110  00001");
    apply_vector ( 9'b100011110,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 100010001  10001");
    apply_vector ( 9'b100010001,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 100011001  01001");
    apply_vector ( 9'b100011001,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 100010101  11001");
    apply_vector ( 9'b100010101,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 100011101  00101");
    apply_vector ( 9'b100011101,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 100010011  10101");
    apply_vector ( 9'b100010011,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 100011011  01101");
    apply_vector ( 9'b100011011,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 100010111  11101");
    apply_vector ( 9'b100010111,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 100011111  00011");
    apply_vector ( 9'b100011111,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 110010000  01010");
    apply_vector ( 9'b110010000,5'b01010,
                   9'b111111111,5'b11111);
    $display ( "v 110011000  11010");
    apply_vector ( 9'b110011000,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 110010100  00110");
    apply_vector ( 9'b110010100,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 110011100  10110");
    apply_vector ( 9'b110011100,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 110010010  01110");
    apply_vector ( 9'b110010010,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 110011010  11110");
    apply_vector ( 9'b110011010,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 110010110  00001");
    apply_vector ( 9'b110010110,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 110011110  10001");
    apply_vector ( 9'b110011110,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 110010001  01001");
    apply_vector ( 9'b110010001,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 110011001  11001");
    apply_vector ( 9'b110011001,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 110010101  00101");
    apply_vector ( 9'b110010101,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 110011101  10101");
    apply_vector ( 9'b110011101,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 110010011  01101");
    apply_vector ( 9'b110010011,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 110011011  11101");
    apply_vector ( 9'b110011011,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 110010111  00011");
    apply_vector ( 9'b110010111,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 110011111  10011");
    apply_vector ( 9'b110011111,5'b10011,
                   9'b111111111,5'b11111);
    $display ( "v 101010000  11010");
    apply_vector ( 9'b101010000,5'b11010,
                   9'b111111111,5'b11111);
    $display ( "v 101011000  00110");
    apply_vector ( 9'b101011000,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 101010100  10110");
    apply_vector ( 9'b101010100,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 101011100  01110");
    apply_vector ( 9'b101011100,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 101010010  11110");
    apply_vector ( 9'b101010010,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 101011010  00001");
    apply_vector ( 9'b101011010,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 101010110  10001");
    apply_vector ( 9'b101010110,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 101011110  01001");
    apply_vector ( 9'b101011110,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 101010001  11001");
    apply_vector ( 9'b101010001,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 101011001  00101");
    apply_vector ( 9'b101011001,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 101010101  10101");
    apply_vector ( 9'b101010101,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 101011101  01101");
    apply_vector ( 9'b101011101,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 101010011  11101");
    apply_vector ( 9'b101010011,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 101011011  00011");
    apply_vector ( 9'b101011011,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 101010111  10011");
    apply_vector ( 9'b101010111,5'b10011,
                   9'b111111111,5'b11111);
    $display ( "v 101011111  01011");
    apply_vector ( 9'b101011111,5'b01011,
                   9'b111111111,5'b11111);
    $display ( "v 111010000  00110");
    apply_vector ( 9'b111010000,5'b00110,
                   9'b111111111,5'b11111);
    $display ( "v 111011000  10110");
    apply_vector ( 9'b111011000,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 111010100  01110");
    apply_vector ( 9'b111010100,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 111011100  11110");
    apply_vector ( 9'b111011100,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 111010010  00001");
    apply_vector ( 9'b111010010,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 111011010  10001");
    apply_vector ( 9'b111011010,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 111010110  01001");
    apply_vector ( 9'b111010110,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 111011110  11001");
    apply_vector ( 9'b111011110,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 111010001  00101");
    apply_vector ( 9'b111010001,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 111011001  10101");
    apply_vector ( 9'b111011001,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 111010101  01101");
    apply_vector ( 9'b111010101,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 111011101  11101");
    apply_vector ( 9'b111011101,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 111010011  00011");
    apply_vector ( 9'b111010011,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 111011011  10011");
    apply_vector ( 9'b111011011,5'b10011,
                   9'b111111111,5'b11111);
    $display ( "v 111010111  01011");
    apply_vector ( 9'b111010111,5'b01011,
                   9'b111111111,5'b11111);
    $display ( "v 111011111  11011");
    apply_vector ( 9'b111011111,5'b11011,
                   9'b111111111,5'b11111);
    $display ( "v 100110000  10110");
    apply_vector ( 9'b100110000,5'b10110,
                   9'b111111111,5'b11111);
    $display ( "v 100111000  01110");
    apply_vector ( 9'b100111000,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 100110100  11110");
    apply_vector ( 9'b100110100,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 100111100  00001");
    apply_vector ( 9'b100111100,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 100110010  10001");
    apply_vector ( 9'b100110010,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 100111010  01001");
    apply_vector ( 9'b100111010,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 100110110  11001");
    apply_vector ( 9'b100110110,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 100111110  00101");
    apply_vector ( 9'b100111110,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 100110001  10101");
    apply_vector ( 9'b100110001,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 100111001  01101");
    apply_vector ( 9'b100111001,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 100110101  11101");
    apply_vector ( 9'b100110101,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 100111101  00011");
    apply_vector ( 9'b100111101,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 100110011  10011");
    apply_vector ( 9'b100110011,5'b10011,
                   9'b111111111,5'b11111);
    $display ( "v 100111011  01011");
    apply_vector ( 9'b100111011,5'b01011,
                   9'b111111111,5'b11111);
    $display ( "v 100110111  11011");
    apply_vector ( 9'b100110111,5'b11011,
                   9'b111111111,5'b11111);
    $display ( "v 100111111  00111");
    apply_vector ( 9'b100111111,5'b00111,
                   9'b111111111,5'b11111);
    $display ( "v 110110000  01110");
    apply_vector ( 9'b110110000,5'b01110,
                   9'b111111111,5'b11111);
    $display ( "v 110111000  11110");
    apply_vector ( 9'b110111000,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 110110100  00001");
    apply_vector ( 9'b110110100,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 110111100  10001");
    apply_vector ( 9'b110111100,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 110110010  01001");
    apply_vector ( 9'b110110010,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 110111010  11001");
    apply_vector ( 9'b110111010,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 110110110  00101");
    apply_vector ( 9'b110110110,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 110111110  10101");
    apply_vector ( 9'b110111110,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 110110001  01101");
    apply_vector ( 9'b110110001,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 110111001  11101");
    apply_vector ( 9'b110111001,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 110110101  00011");
    apply_vector ( 9'b110110101,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 110111101  10011");
    apply_vector ( 9'b110111101,5'b10011,
                   9'b111111111,5'b11111);
    $display ( "v 110110011  01011");
    apply_vector ( 9'b110110011,5'b01011,
                   9'b111111111,5'b11111);
    $display ( "v 110111011  11011");
    apply_vector ( 9'b110111011,5'b11011,
                   9'b111111111,5'b11111);
    $display ( "v 110110111  00111");
    apply_vector ( 9'b110110111,5'b00111,
                   9'b111111111,5'b11111);
    $display ( "v 110111111  10111");
    apply_vector ( 9'b110111111,5'b10111,
                   9'b111111111,5'b11111);
    $display ( "v 101110000  11110");
    apply_vector ( 9'b101110000,5'b11110,
                   9'b111111111,5'b11111);
    $display ( "v 101111000  00001");
    apply_vector ( 9'b101111000,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 101110100  10001");
    apply_vector ( 9'b101110100,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 101111100  01001");
    apply_vector ( 9'b101111100,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 101110010  11001");
    apply_vector ( 9'b101110010,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 101111010  00101");
    apply_vector ( 9'b101111010,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 101110110  10101");
    apply_vector ( 9'b101110110,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 101111110  01101");
    apply_vector ( 9'b101111110,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 101110001  11101");
    apply_vector ( 9'b101110001,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 101111001  00011");
    apply_vector ( 9'b101111001,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 101110101  10011");
    apply_vector ( 9'b101110101,5'b10011,
                   9'b111111111,5'b11111);
    $display ( "v 101111101  01011");
    apply_vector ( 9'b101111101,5'b01011,
                   9'b111111111,5'b11111);
    $display ( "v 101110011  11011");
    apply_vector ( 9'b101110011,5'b11011,
                   9'b111111111,5'b11111);
    $display ( "v 101111011  00111");
    apply_vector ( 9'b101111011,5'b00111,
                   9'b111111111,5'b11111);
    $display ( "v 101110111  10111");
    apply_vector ( 9'b101110111,5'b10111,
                   9'b111111111,5'b11111);
    $display ( "v 101111111  01111");
    apply_vector ( 9'b101111111,5'b01111,
                   9'b111111111,5'b11111);
    $display ( "v 111110000  00001");
    apply_vector ( 9'b111110000,5'b00001,
                   9'b111111111,5'b11111);
    $display ( "v 111111000  10001");
    apply_vector ( 9'b111111000,5'b10001,
                   9'b111111111,5'b11111);
    $display ( "v 111110100  01001");
    apply_vector ( 9'b111110100,5'b01001,
                   9'b111111111,5'b11111);
    $display ( "v 111111100  11001");
    apply_vector ( 9'b111111100,5'b11001,
                   9'b111111111,5'b11111);
    $display ( "v 111110010  00101");
    apply_vector ( 9'b111110010,5'b00101,
                   9'b111111111,5'b11111);
    $display ( "v 111111010  10101");
    apply_vector ( 9'b111111010,5'b10101,
                   9'b111111111,5'b11111);
    $display ( "v 111110110  01101");
    apply_vector ( 9'b111110110,5'b01101,
                   9'b111111111,5'b11111);
    $display ( "v 111111110  11101");
    apply_vector ( 9'b111111110,5'b11101,
                   9'b111111111,5'b11111);
    $display ( "v 111110001  00011");
    apply_vector ( 9'b111110001,5'b00011,
                   9'b111111111,5'b11111);
    $display ( "v 111111001  10011");
    apply_vector ( 9'b111111001,5'b10011,
                   9'b111111111,5'b11111);
    $display ( "v 111110101  01011");
    apply_vector ( 9'b111110101,5'b01011,
                   9'b111111111,5'b11111);
    $display ( "v 111111101  11011");
    apply_vector ( 9'b111111101,5'b11011,
                   9'b111111111,5'b11111);
    $display ( "v 111110011  00111");
    apply_vector ( 9'b111110011,5'b00111,
                   9'b111111111,5'b11111);
    $display ( "v 111111011  10111");
    apply_vector ( 9'b111111011,5'b10111,
                   9'b111111111,5'b11111);
    $display ( "v 111110111  01111");
    apply_vector ( 9'b111110111,5'b01111,
                   9'b111111111,5'b11111);
    $display ( "v 111111111  11111");
    apply_vector ( 9'b111111111,5'b11111,
                   9'b111111111,5'b11111);
    if ( errors == 0 )
      begin
        $display( "Simulation OK" );
        $display( "All vectors passed" );
      end
    else
      begin
        $display( "" );
        $display( "Simulation Failed" );
        $display( "" );
        if (  errors_Q3 > 0 )
          $display ( "       ", errors_Q3, " errors with Q3",) ;
        if (  errors_Q4 > 0 )
          $display ( "       ", errors_Q4, " errors with Q4",) ;
        if (  errors_Q5 > 0 )
          $display ( "       ", errors_Q5, " errors with Q5",) ;
        if (  errors_Q6 > 0 )
          $display ( "       ", errors_Q6, " errors with Q6",) ;
        if (  errors_Q7 > 0 )
          $display ( "       ", errors_Q7, " errors with Q7",) ;
        $display( "" );
        $display( "Total: ", errors, " errors");
        $display( "" );
      end
    $stop;
    $finish;
  end

// function declaration

task apply_vector;

  input [8:0] stimulus_vector;
  input [4:0] expected_vector;
  input [8:0] stimulus_mask;
  input [4:0] expected_mask;

  begin
    `ifdef set_x_to_0
      {A3,A4,A5,A6,A7,A8,A9,A10,A11} = stimulus_vector & stimulus_mask ;
    `else
      {A3,A4,A5,A6,A7,A8,A9,A10,A11} = stimulus_vector;
    `endif
    #500
    check_vector( expected_vector, expected_mask );
    #500
    $display("");
  end

endtask
task check_vector;

  input [4:0] expected_vector;
  input [4:0] mask_vector;

  reg [4:0] received_vector;
  reg [4:0] difference_vector;

  integer local_errors;

  begin
    local_errors = 0;
    received_vector = {Q3,Q4,Q5,Q6,Q7};
    difference_vector = ( received_vector ^ expected_vector ) & mask_vector ;
    $display( "r            %b", received_vector );
    $display( "             %s", error_point( difference_vector ) );
    if ( expected_vector[4] !== 1'bX )
      if ( expected_vector[4] !== Q3)
        begin
          $display( "error with Q3 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q3 = errors_Q3 + 1;
        end
    if ( expected_vector[3] !== 1'bX )
      if ( expected_vector[3] !== Q4)
        begin
          $display( "error with Q4 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q4 = errors_Q4 + 1;
        end
    if ( expected_vector[2] !== 1'bX )
      if ( expected_vector[2] !== Q5)
        begin
          $display( "error with Q5 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q5 = errors_Q5 + 1;
        end
    if ( expected_vector[1] !== 1'bX )
      if ( expected_vector[1] !== Q6)
        begin
          $display( "error with Q6 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q6 = errors_Q6 + 1;
        end
    if ( expected_vector[0] !== 1'bX )
      if ( expected_vector[0] !== Q7)
        begin
          $display( "error with Q7 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q7 = errors_Q7 + 1;
        end
    if ( local_errors > 0 ) $display( "" );
    errors = errors + local_errors;
  end

endtask
function [39:0] error_point;

  input [4:0] in_vector;
  integer i, j;
  begin
    error_point[ 7 : 0 ] = ( in_vector[ 0 ] === 0 ) ? " " : "^";
    error_point[ 15 : 8 ] = ( in_vector[ 1 ] === 0 ) ? " " : "^";
    error_point[ 23 : 16 ] = ( in_vector[ 2 ] === 0 ) ? " " : "^";
    error_point[ 31 : 24 ] = ( in_vector[ 3 ] === 0 ) ? " " : "^";
    error_point[ 39 : 32 ] = ( in_vector[ 4 ] === 0 ) ? " " : "^";
  end

endfunction


endmodule

