// Verilog test bench for D2 chip design

`timescale 1ns/1ps

module test_TEAMJ_DESIGN;

// declare DUT input signals as "reg"
// declare DUT output signals as "wire"

reg A0;
reg A1;
reg A2;
reg A3;
reg A4;
reg A5;
reg A6;
reg A7;
reg A8;
reg A9;
reg A10;
reg A11;
reg A12;
reg A13;
reg A14;
reg A15;
reg A16;
reg A17;
reg A18;
reg A19;
reg A20;
reg A21;
reg A22;
reg A23;
wire Q0;
wire Q1;
wire Q3;
wire Q4;
wire Q5;
wire Q6;
wire Q7;
wire Q12;
wire Q15;
wire Q16;
wire Q17;
wire Q18;
wire Q19;
wire Q20;
wire Q21;
wire Q22;
wire Q23;
integer errors_Q0;
integer errors_Q1;
integer errors_Q3;
integer errors_Q4;
integer errors_Q5;
integer errors_Q6;
integer errors_Q7;
integer errors_Q12;
integer errors_Q15;
integer errors_Q16;
integer errors_Q17;
integer errors_Q18;
integer errors_Q19;
integer errors_Q20;
integer errors_Q21;
integer errors_Q22;
integer errors_Q23;

// declare error count

integer errors;

// instance Device Under Test
//   assumes top-level OrCAD schematic is named "TEAMJ_DESIGN"

`ifdef DUT
  `DUT DUT(
`else
  TEAMJ_DESIGN DUT(
`endif
   .A0(A0),
   .A1(A1),
   .A2(A2),
   .A3(A3),
   .A4(A4),
   .A5(A5),
   .A6(A6),
   .A7(A7),
   .A8(A8),
   .A9(A9),
   .A10(A10),
   .A11(A11),
   .A12(A12),
   .A13(A13),
   .A14(A14),
   .A15(A15),
   .A16(A16),
   .A17(A17),
   .A18(A18),
   .A19(A19),
   .A20(A20),
   .A21(A21),
   .A22(A22),
   .A23(A23),
   .Q0(Q0),
   .Q1(Q1),
   .Q3(Q3),
   .Q4(Q4),
   .Q5(Q5),
   .Q6(Q6),
   .Q7(Q7),
   .Q12(Q12),
   .Q15(Q15),
   .Q16(Q16),
   .Q17(Q17),
   .Q18(Q18),
   .Q19(Q19),
   .Q20(Q20),
   .Q21(Q21),
   .Q22(Q22),
   .Q23(Q23)
);

// monitor the I/O
initial
  begin
    $display( "Simulation Begins" );
    $display ( "  AAAAAAAAAAAAAAAAAAAAAAAA  QQQQQQQQQQQQQQQQQ" );
    $display ( "  012345678911111111112222  01345671111112222" );
    $display ( "            01234567890123         2567890123" );
    $display ( "                                             " );
    `ifdef no_monitor
    `else
    $monitor ( "  ",
      A0,
      A1,
      A2,
      A3,
      A4,
      A5,
      A6,
      A7,
      A8,
      A9,
      A10,
      A11,
      A12,
      A13,
      A14,
      A15,
      A16,
      A17,
      A18,
      A19,
      A20,
      A21,
      A22,
      A23,
      "  ",
      Q0,
      Q1,
      Q3,
      Q4,
      Q5,
      Q6,
      Q7,
      Q12,
      Q15,
      Q16,
      Q17,
      Q18,
      Q19,
      Q20,
      Q21,
      Q22,
      Q23,
      "  @ %d ns", $time   );
    `endif
  end

// stimulii

initial
  begin
    errors = 0;
    errors_Q0 = 0;
    errors_Q1 = 0;
    errors_Q3 = 0;
    errors_Q4 = 0;
    errors_Q5 = 0;
    errors_Q6 = 0;
    errors_Q7 = 0;
    errors_Q12 = 0;
    errors_Q15 = 0;
    errors_Q16 = 0;
    errors_Q17 = 0;
    errors_Q18 = 0;
    errors_Q19 = 0;
    errors_Q20 = 0;
    errors_Q21 = 0;
    errors_Q22 = 0;
    errors_Q23 = 0;
    $display ( "v 001000000000000000000000  10000000000000000");
    apply_vector ( 24'b001000000000000000000000,17'b10000000000000000,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111000001000000000000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000000000000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000000100000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000000100000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000000000000000  0X100000000000000");
    apply_vector ( 24'b111000001000000000000000,17'b0X100000000000000,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010000000100000011000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100000011000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100000111000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100000111000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100000011000010  11010000110000000");
    apply_vector ( 24'b010000000100000011000010,17'b11010000110000000,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111000001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100000010000000  0X110000000000000");
    apply_vector ( 24'b111000001100000010000000,17'b0X110000000000000,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001000000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010000010000000  10001000010000000");
    apply_vector ( 24'b001000000010000010000000,17'b10001000010000000,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111000001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010000010000000  0X101000000000000");
    apply_vector ( 24'b111000001010000010000000,17'b0X101000000000000,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010000000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110000010000000  11011000010000000");
    apply_vector ( 24'b010000000110000010000000,17'b11011000010000000,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111000001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110000010000000  0X111000000000000");
    apply_vector ( 24'b111000001110000010000000,17'b0X111000000000000,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001000000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001000010000000  10000100000000000");
    apply_vector ( 24'b001000000001000010000000,17'b10000100000000000,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111000001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001000010000000  0X100100001100011");
    apply_vector ( 24'b111000001001000010000000,17'b0X100100001100011,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010000000101000011100011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101000011100011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101000111100011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101000111100011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101000011100011  11010100100100010");
    apply_vector ( 24'b010000000101000011100011,17'b11010100100100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111000001101000010100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101000010100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101000110100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101000110100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101000010100000  0X110100010100010");
    apply_vector ( 24'b111000001101000010100000,17'b0X110100010100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001000000011000010100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011000010100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011000110100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011000110100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011000010100000  10001100000100010");
    apply_vector ( 24'b001000000011000010100000,17'b10001100000100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111000001011000010100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011000010100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011000110100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011000110100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011000010100000  0X101100000100010");
    apply_vector ( 24'b111000001011000010100000,17'b0X101100000100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010000000111000010100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111000010100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111000110100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111000110100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111000010100000  11011100000100010");
    apply_vector ( 24'b010000000111000010100000,17'b11011100000100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111000001111000010100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111000010100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111000110100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111000110100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111000010100000  0X111100000100010");
    apply_vector ( 24'b111000001111000010100000,17'b0X111100000100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001010000000000010100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000000010100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000000110100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000000110100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000000010100000  10100000000100010");
    apply_vector ( 24'b001010000000000010100000,17'b10100000000100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111010001000000010100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000000010100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000000110100000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000000110100000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000000010100000  0X010000001XXXX01");
    apply_vector ( 24'b111010001000000010100000,17'b0X010000001XXXX01,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010010000100000011010010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100000011010010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100000111010010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100000111010010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100000011010010  11110000110XXXX00");
    apply_vector ( 24'b010010000100000011010010,17'b11110000110XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111010001100000010010001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100000010010001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100000110010001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100000110010001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100000010010001  0X001000000XXXX00");
    apply_vector ( 24'b111010001100000010010001,17'b0X001000000XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001010000010000010010000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010000010010000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010000110010000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010000110010000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010000010010000  10101000000XXXX00");
    apply_vector ( 24'b001010000010000010010000,17'b10101000000XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111010001010000010010000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010000010010000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010000110010000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010000110010000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010000010010000  0X011000010XXXX00");
    apply_vector ( 24'b111010001010000010010000,17'b0X011000010XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010010000110000010010000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110000010010000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110000110010000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110000110010000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110000010010000  11111000000XXXX00");
    apply_vector ( 24'b010010000110000010010000,17'b11111000000XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111010001110000010010000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110000010010000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110000110010000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110000110010000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110000010010000  0X000100000XXXX00");
    apply_vector ( 24'b111010001110000010010000,17'b0X000100000XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001010000001000010010000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001000010010000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001000110010000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001000110010000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001000010010000  10100100010XXXX00");
    apply_vector ( 24'b001010000001000010010000,17'b10100100010XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111010001001000010010000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001000010010000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001000110010000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001000110010000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001000010010000  0X010100001100010");
    apply_vector ( 24'b111010001001000010010000,17'b0X010100001100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010010000101000011110011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101000011110011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101000111110011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101000111110011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101000011110011  11110100100100010");
    apply_vector ( 24'b010010000101000011110011,17'b11110100100100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111010001101000010110001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101000010110001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101000110110001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101000110110001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101000010110001  0X001100010100010");
    apply_vector ( 24'b111010001101000010110001,17'b0X001100010100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001010000011000010110000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011000010110000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011000110110000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011000110110000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011000010110000  10101100010100010");
    apply_vector ( 24'b001010000011000010110000,17'b10101100010100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111010001011000010110000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011000010110000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011000110110000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011000110110000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011000010110000  0X011100010100010");
    apply_vector ( 24'b111010001011000010110000,17'b0X011100010100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010010000111000010110000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111000010110000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111000110110000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111000110110000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111000010110000  11111100010100010");
    apply_vector ( 24'b010010000111000010110000,17'b11111100010100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111010001111000010110000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111000010110000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111000110110000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111000110110000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111000010110000  0X000010000100010");
    apply_vector ( 24'b111010001111000010110000,17'b0X000010000100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001001000000000010110000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000000010110000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000000110110000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000000110110000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000000010110000  10010000010100010");
    apply_vector ( 24'b001001000000000010110000,17'b10010000010100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111001001000000010110000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000000010110000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000000110110000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000000110110000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000000010110000  0X110000001100011");
    apply_vector ( 24'b111001001000000010110000,17'b0X110000001100011,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010001000100000011001010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100000011001010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100000111001010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100000111001010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100000011001010  11001000100100010");
    apply_vector ( 24'b010001000100000011001010,17'b11001000100100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111001001100000010001000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100000010001000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100000110001000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100000110001000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100000010001000  0X101000000100010");
    apply_vector ( 24'b111001001100000010001000,17'b0X101000000100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001001000010000010001001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010000010001001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010000110001001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010000110001001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010000010001001  10011000010100010");
    apply_vector ( 24'b001001000010000010001001,17'b10011000010100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111001001010000010001000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010000010001000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010000110001000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010000110001000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010000010001000  0X111000000100010");
    apply_vector ( 24'b111001001010000010001000,17'b0X111000000100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010001000110000010001000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110000010001000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110000110001000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110000110001000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110000010001000  11000100000100010");
    apply_vector ( 24'b010001000110000010001000,17'b11000100000100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111001001110000010001000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110000010001000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110000110001000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110000110001000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110000010001000  0X100100010100010");
    apply_vector ( 24'b111001001110000010001000,17'b0X100100010100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001001000001000010001000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001000010001000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001000110001000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001000110001000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001000010001000  10010100010100010");
    apply_vector ( 24'b001001000001000010001000,17'b10010100010100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111001001001000010001000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001000010001000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001000110001000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001000110001000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001000010001000  0X110100001XXXX01");
    apply_vector ( 24'b111001001001000010001000,17'b0X110100001XXXX01,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010001000101000011101011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101000011101011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101000111101011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101000111101011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101000011101011  11001100110XXXX00");
    apply_vector ( 24'b010001000101000011101011,17'b11001100110XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111001001101000010101000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101000010101000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101000110101000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101000110101000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101000010101000  0X101100010XXXX00");
    apply_vector ( 24'b111001001101000010101000,17'b0X101100010XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001001000011000010101001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011000010101001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011000110101001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011000110101001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011000010101001  10011100000XXXX00");
    apply_vector ( 24'b001001000011000010101001,17'b10011100000XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111001001011000010101000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011000010101000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011000110101000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011000110101000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011000010101000  0X111100000XXXX00");
    apply_vector ( 24'b111001001011000010101000,17'b0X111100000XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010001000111000010101000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111000010101000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111000110101000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111000110101000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111000010101000  11000010010XXXX00");
    apply_vector ( 24'b010001000111000010101000,17'b11000010010XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111001001111000010101000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111000010101000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111000110101000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111000110101000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111000010101000  0X100010010XXXX00");
    apply_vector ( 24'b111001001111000010101000,17'b0X100010010XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001011000000000010101000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000000010101000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000000110101000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000000110101000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000000010101000  10110000010XXXX00");
    apply_vector ( 24'b001011000000000010101000,17'b10110000010XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111011001000000010101000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000000010101000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000000110101000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000000110101000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000000010101000  0X001000001000011");
    apply_vector ( 24'b111011001000000010101000,17'b0X001000001000011,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010011000100000011011010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100000011011010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100000111011010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100000111011010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100000011011010  11101000100000010");
    apply_vector ( 24'b010011000100000011011010,17'b11101000100000010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111011001100000010011001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100000010011001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100000110011001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100000110011001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100000010011001  0X011000000000010");
    apply_vector ( 24'b111011001100000010011001,17'b0X011000000000010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001011000010000010011001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010000010011001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010000110011001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010000110011001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010000010011001  10111000000000010");
    apply_vector ( 24'b001011000010000010011001,17'b10111000000000010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111011001010000010011000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010000010011000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010000110011000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010000110011000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010000010011000  0X000100010000010");
    apply_vector ( 24'b111011001010000010011000,17'b0X000100010000010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010011000110000010011000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110000010011000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110000110011000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110000110011000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110000010011000  11100100010000010");
    apply_vector ( 24'b010011000110000010011000,17'b11100100010000010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111011001110000010011000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110000010011000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110000110011000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110000110011000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110000010011000  0X010100010000010");
    apply_vector ( 24'b111011001110000010011000,17'b0X010100010000010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001011000001000010011000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001000010011000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001000110011000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001000110011000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001000010011000  10110100000000010");
    apply_vector ( 24'b001011000001000010011000,17'b10110100000000010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111011001001000010011000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001000010011000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001000110011000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001000110011000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001000010011000  0X001100001100011");
    apply_vector ( 24'b111011001001000010011000,17'b0X001100001100011,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010011000101000011111011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101000011111011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101000111111011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101000111111011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101000011111011  11101100110100010");
    apply_vector ( 24'b010011000101000011111011,17'b11101100110100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111011001101000010111001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101000010111001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101000110111001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101000110111001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101000010111001  0X011100010100010");
    apply_vector ( 24'b111011001101000010111001,17'b0X011100010100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001011000011000010111001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011000010111001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011000110111001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011000110111001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011000010111001  10111100010100010");
    apply_vector ( 24'b001011000011000010111001,17'b10111100010100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111011001011000010111000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011000010111000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011000110111000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011000110111000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011000010111000  0X000010010100010");
    apply_vector ( 24'b111011001011000010111000,17'b0X000010010100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010011000111000010111000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111000010111000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111000110111000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111000110111000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111000010111000  11100010000100010");
    apply_vector ( 24'b010011000111000010111000,17'b11100010000100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111011001111000010111000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111000010111000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111000110111000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111000110111000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111000010111000  0X010010010100010");
    apply_vector ( 24'b111011001111000010111000,17'b0X010010010100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001000100000000010111000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000000010111000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000000110111000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000000110111000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000000010111000  10001000000100010");
    apply_vector ( 24'b001000100000000010111000,17'b10001000000100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111000101000000010111000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000000010111000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000000110111000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000000110111000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000000010111000  0X101000001XXXX01");
    apply_vector ( 24'b111000101000000010111000,17'b0X101000001XXXX01,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010000100100000011000110  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100000011000110,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100000111000110  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100000111000110,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100000011000110  11011000100XXXX00");
    apply_vector ( 24'b010000100100000011000110,17'b11011000100XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111000101100000010000100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100000010000100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100000110000100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100000110000100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100000010000100  0X111000000XXXX00");
    apply_vector ( 24'b111000101100000010000100,17'b0X111000000XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001000100010000010000100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010000010000100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010000110000100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010000110000100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010000010000100  10000100000XXXX00");
    apply_vector ( 24'b001000100010000010000100,17'b10000100000XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111000101010000010000101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010000010000101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010000110000101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010000110000101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010000010000101  0X100100000XXXX00");
    apply_vector ( 24'b111000101010000010000101,17'b0X100100000XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010000100110000010000100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110000010000100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110000110000100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110000110000100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110000010000100  11010100010XXXX00");
    apply_vector ( 24'b010000100110000010000100,17'b11010100010XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111000101110000010000100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110000010000100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110000110000100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110000110000100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110000010000100  0X110100000XXXX00");
    apply_vector ( 24'b111000101110000010000100,17'b0X110100000XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001000100001000010000100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001000010000100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001000110000100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001000110000100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001000010000100  10001100010XXXX00");
    apply_vector ( 24'b001000100001000010000100,17'b10001100010XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111000101001000010000100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001000010000100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001000110000100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001000110000100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001000010000100  0X101100011XXXX01");
    apply_vector ( 24'b111000101001000010000100,17'b0X101100011XXXX01,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010000100101000011100111  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101000011100111,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101000111100111  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101000111100111,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101000011100111  11011100110XXXX00");
    apply_vector ( 24'b010000100101000011100111,17'b11011100110XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111000101101000010100100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101000010100100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101000110100100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101000110100100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101000010100100  0X111100010XXXX00");
    apply_vector ( 24'b111000101101000010100100,17'b0X111100010XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001000100011000010100100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011000010100100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011000110100100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011000110100100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011000010100100  10000010010XXXX00");
    apply_vector ( 24'b001000100011000010100100,17'b10000010010XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111000101011000010100101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011000010100101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011000110100101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011000110100101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011000010100101  0X100010000XXXX00");
    apply_vector ( 24'b111000101011000010100101,17'b0X100010000XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010000100111000010100100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111000010100100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111000110100100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111000110100100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111000010100100  11010010000XXXX00");
    apply_vector ( 24'b010000100111000010100100,17'b11010010000XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111000101111000010100100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111000010100100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111000110100100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111000110100100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111000010100100  0X110010000XXXX00");
    apply_vector ( 24'b111000101111000010100100,17'b0X110010000XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001010100000000010100100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000000010100100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000000110100100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000000110100100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000000010100100  10101000010XXXX00");
    apply_vector ( 24'b001010100000000010100100,17'b10101000010XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111010101000000010100100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000000010100100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000000110100100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000000110100100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000000010100100  0X011000011010011");
    apply_vector ( 24'b111010101000000010100100,17'b0X011000011010011,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010010100100000011010110  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100000011010110,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100000111010110  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100000111010110,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100000011010110  11111000100010010");
    apply_vector ( 24'b010010100100000011010110,17'b11111000100010010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111010101100000010010101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100000010010101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100000110010101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100000110010101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100000010010101  0X000100000010010");
    apply_vector ( 24'b111010101100000010010101,17'b0X000100000010010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001010100010000010010100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010000010010100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010000110010100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010000110010100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010000010010100  10100100010010010");
    apply_vector ( 24'b001010100010000010010100,17'b10100100010010010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111010101010000010010101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010000010010101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010000110010101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010000110010101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010000010010101  0X010100010010010");
    apply_vector ( 24'b111010101010000010010101,17'b0X010100010010010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010010100110000010010100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110000010010100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110000110010100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110000110010100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110000010010100  11110100000010010");
    apply_vector ( 24'b010010100110000010010100,17'b11110100000010010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111010101110000010010100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110000010010100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110000110010100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110000110010100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110000010010100  0X001100000010010");
    apply_vector ( 24'b111010101110000010010100,17'b0X001100000010010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001010100001000010010100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001000010010100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001000110010100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001000110010100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001000010010100  10101100000010010");
    apply_vector ( 24'b001010100001000010010100,17'b10101100000010010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111010101001000010010100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001000010010100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001000110010100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001000110010100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001000010010100  0X011100011100011");
    apply_vector ( 24'b111010101001000010010100,17'b0X011100011100011,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010010100101000011110111  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101000011110111,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101000111110111  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101000111110111,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101000011110111  11111100110100010");
    apply_vector ( 24'b010010100101000011110111,17'b11111100110100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111010101101000010110101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101000010110101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101000110110101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101000110110101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101000010110101  0X000010010100010");
    apply_vector ( 24'b111010101101000010110101,17'b0X000010010100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001010100011000010110100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011000010110100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011000110110100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011000110110100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011000010110100  10100010000100010");
    apply_vector ( 24'b001010100011000010110100,17'b10100010000100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111010101011000010110101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011000010110101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011000110110101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011000110110101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011000010110101  0X010010010100010");
    apply_vector ( 24'b111010101011000010110101,17'b0X010010010100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010010100111000010110100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111000010110100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111000110110100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111000110110100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111000010110100  11110010010100010");
    apply_vector ( 24'b010010100111000010110100,17'b11110010010100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111010101111000010110100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111000010110100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111000110110100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111000110110100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111000010110100  0X001010000100010");
    apply_vector ( 24'b111010101111000010110100,17'b0X001010000100010,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001001100000000010110100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000000010110100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000000110110100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000000110110100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000000010110100  10011000000100010");
    apply_vector ( 24'b001001100000000010110100,17'b10011000000100010,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111001101000000010110100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000000010110100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000000110110100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000000110110100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000000010110100  0X111000011XXXX01");
    apply_vector ( 24'b111001101000000010110100,17'b0X111000011XXXX01,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010001100100000011001110  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100000011001110,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100000111001110  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100000111001110,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100000011001110  11000100110XXXX00");
    apply_vector ( 24'b010001100100000011001110,17'b11000100110XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111001101100000010001100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100000010001100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100000110001100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100000110001100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100000010001100  0X100100000XXXX00");
    apply_vector ( 24'b111001101100000010001100,17'b0X100100000XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001001100010000010001101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010000010001101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010000110001101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010000110001101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010000010001101  10010100000XXXX00");
    apply_vector ( 24'b001001100010000010001101,17'b10010100000XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111001101010000010001101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010000010001101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010000110001101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010000110001101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010000010001101  0X110100000XXXX00");
    apply_vector ( 24'b111001101010000010001101,17'b0X110100000XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010001100110000010001100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110000010001100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110000110001100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110000110001100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110000010001100  11001100000XXXX00");
    apply_vector ( 24'b010001100110000010001100,17'b11001100000XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111001101110000010001100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110000010001100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110000110001100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110000110001100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110000010001100  0X101100010XXXX00");
    apply_vector ( 24'b111001101110000010001100,17'b0X101100010XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001001100001000010001100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001000010001100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001000110001100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001000110001100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001000010001100  10011100000XXXX00");
    apply_vector ( 24'b001001100001000010001100,17'b10011100000XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111001101001000010001100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001000010001100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001000110001100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001000110001100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001000010001100  0X111100011010111");
    apply_vector ( 24'b111001101001000010001100,17'b0X111100011010111,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010001100101000011101111  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101000011101111,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101000111101111  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101000111101111,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101000011101111  11000010100010110");
    apply_vector ( 24'b010001100101000011101111,17'b11000010100010110,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111001101101000010101100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101000010101100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101000110101100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101000110101100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101000010101100  0X100010010010110");
    apply_vector ( 24'b111001101101000010101100,17'b0X100010010010110,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001001100011000010101101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011000010101101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011000110101101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011000110101101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011000010101101  10010010010010110");
    apply_vector ( 24'b001001100011000010101101,17'b10010010010010110,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111001101011000010101101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011000010101101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011000110101101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011000110101101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011000010101101  0X110010000010110");
    apply_vector ( 24'b111001101011000010101101,17'b0X110010000010110,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010001100111000010101100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111000010101100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111000110101100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111000110101100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111000010101100  11001010010010110");
    apply_vector ( 24'b010001100111000010101100,17'b11001010010010110,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111001101111000010101100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111000010101100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111000110101100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111000110101100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111000010101100  0X101010010010110");
    apply_vector ( 24'b111001101111000010101100,17'b0X101010010010110,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 001011100000000010101100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000000010101100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000000110101100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000000110101100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000000010101100  10111000000010110");
    apply_vector ( 24'b001011100000000010101100,17'b10111000000010110,
                   24'b111111111111111111111111,17'b11111111111111111);
    $display ( "v 111011101000000010101100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000000010101100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000000110101100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000000110101100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000000010101100  0X000100011XXXX01");
    apply_vector ( 24'b111011101000000010101100,17'b0X000100011XXXX01,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010011100100000011011110  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100000011011110,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100000111011110  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100000111011110,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100000011011110  11100100110XXXX00");
    apply_vector ( 24'b010011100100000011011110,17'b11100100110XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111011101100000010011101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100000010011101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100000110011101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100000110011101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100000010011101  0X010100000XXXX00");
    apply_vector ( 24'b111011101100000010011101,17'b0X010100000XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001011100010000010011101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010000010011101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010000110011101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010000110011101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010000010011101  10110100010XXXX00");
    apply_vector ( 24'b001011100010000010011101,17'b10110100010XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111011101010000010011101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010000010011101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010000110011101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010000110011101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010000010011101  0X001100010XXXX00");
    apply_vector ( 24'b111011101010000010011101,17'b0X001100010XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010011100110000010011100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110000010011100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110000110011100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110000110011100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110000010011100  11101100010XXXX00");
    apply_vector ( 24'b010011100110000010011100,17'b11101100010XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111011101110000010011100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110000010011100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110000110011100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110000110011100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110000010011100  0X011100010XXXX00");
    apply_vector ( 24'b111011101110000010011100,17'b0X011100010XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001011100001000010011100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001000010011100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001000110011100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001000110011100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001000010011100  10111100010XXXX00");
    apply_vector ( 24'b001011100001000010011100,17'b10111100010XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111011101001000010011100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001000010011100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001000110011100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001000110011100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001000010011100  0X000010011XXXX01");
    apply_vector ( 24'b111011101001000010011100,17'b0X000010011XXXX01,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010011100101000011111111  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101000011111111,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101000111111111  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101000111111111,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101000011111111  11100010100XXXX00");
    apply_vector ( 24'b010011100101000011111111,17'b11100010100XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111011101101000010111101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101000010111101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101000110111101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101000110111101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101000010111101  0X010010010XXXX00");
    apply_vector ( 24'b111011101101000010111101,17'b0X010010010XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001011100011000010111101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011000010111101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011000110111101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011000110111101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011000010111101  10110010000XXXX00");
    apply_vector ( 24'b001011100011000010111101,17'b10110010000XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111011101011000010111101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011000010111101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011000110111101  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011000110111101,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011000010111101  0X001010010XXXX00");
    apply_vector ( 24'b111011101011000010111101,17'b0X001010010XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 010011100111000010111100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111000010111100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111000110111100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111000110111100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111000010111100  11101010000XXXX00");
    apply_vector ( 24'b010011100111000010111100,17'b11101010000XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111011101111000010111100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111000010111100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111000110111100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111000110111100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111000010111100  0X011010010XXXX00");
    apply_vector ( 24'b111011101111000010111100,17'b0X011010010XXXX00,
                   24'b111111111111111111111111,17'b10111111111000011);
    $display ( "v 001000010000000010111100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000000010111100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000000110111100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000000110111100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000000010111100  10000100010XXXX00");
    apply_vector ( 24'b001000010000000010111100,17'b10000100010XXXX00,
                   24'b111111111111111111111111,17'b11111111111000011);
    $display ( "v 111000011000000010111100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000000010111100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000000110111100  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000000110111100,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000000010111100  0X100100011111011");
    apply_vector ( 24'b111000011000000010111100,17'b0X100100011111011,
                   24'b111111111111111111111111,17'b10111111111111111);
    $display ( "v 010000010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100000010000010  110101000X0111010");
    apply_vector ( 24'b010000010100000010000010,17'b110101000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100000010000000  0X1101000X0111010");
    apply_vector ( 24'b111000011100000010000000,17'b0X1101000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010000010000000  100011000X0111010");
    apply_vector ( 24'b001000010010000010000000,17'b100011000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010000010000000  0X1011000X0111010");
    apply_vector ( 24'b111000011010000010000000,17'b0X1011000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110000010000001  110111000X0111010");
    apply_vector ( 24'b010000010110000010000001,17'b110111000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110000010000000  0X1111000X0111010");
    apply_vector ( 24'b111000011110000010000000,17'b0X1111000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001000010000000  100000100X0111010");
    apply_vector ( 24'b001000010001000010000000,17'b100000100X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001000010000000  0X1000100X1XXXX01");
    apply_vector ( 24'b111000011001000010000000,17'b0X1000100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101000010000011  110100100X0XXXX00");
    apply_vector ( 24'b010000010101000010000011,17'b110100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101000010000000  0X1100100X0XXXX00");
    apply_vector ( 24'b111000011101000010000000,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011000010000000  100010100X0XXXX00");
    apply_vector ( 24'b001000010011000010000000,17'b100010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011000010000000  0X1010100X0XXXX00");
    apply_vector ( 24'b111000011011000010000000,17'b0X1010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111000010000001  110110100X0XXXX00");
    apply_vector ( 24'b010000010111000010000001,17'b110110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111000010000000  0X1110100X0XXXX00");
    apply_vector ( 24'b111000011111000010000000,17'b0X1110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000000010000000  101001000X0XXXX00");
    apply_vector ( 24'b001010010000000010000000,17'b101001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000000010000000  0X0101000X1000011");
    apply_vector ( 24'b111010011000000010000000,17'b0X0101000X1000011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100000010000010  111101000X0000010");
    apply_vector ( 24'b010010010100000010000010,17'b111101000X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100000010000001  0X0011000X0000010");
    apply_vector ( 24'b111010011100000010000001,17'b0X0011000X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010000010000000  101011000X0000010");
    apply_vector ( 24'b001010010010000010000000,17'b101011000X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010000010000000  0X0111000X0000010");
    apply_vector ( 24'b111010011010000010000000,17'b0X0111000X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110000010000001  111111000X0000010");
    apply_vector ( 24'b010010010110000010000001,17'b111111000X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110000010000000  0X0000100X0000010");
    apply_vector ( 24'b111010011110000010000000,17'b0X0000100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001000010000000  101000100X0000010");
    apply_vector ( 24'b001010010001000010000000,17'b101000100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001000010000000  0X0100100X1100011");
    apply_vector ( 24'b111010011001000010000000,17'b0X0100100X1100011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101000010000011  111100100X0100010");
    apply_vector ( 24'b010010010101000010000011,17'b111100100X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101000010000001  0X0010100X0100010");
    apply_vector ( 24'b111010011101000010000001,17'b0X0010100X0100010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011000010000000  101010100X0100010");
    apply_vector ( 24'b001010010011000010000000,17'b101010100X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011000010000000  0X0110100X0100010");
    apply_vector ( 24'b111010011011000010000000,17'b0X0110100X0100010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111000010000001  111110100X0100010");
    apply_vector ( 24'b010010010111000010000001,17'b111110100X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111000010000000  0X0001100X0100010");
    apply_vector ( 24'b111010011111000010000000,17'b0X0001100X0100010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000000010000000  100101000X0100010");
    apply_vector ( 24'b001001010000000010000000,17'b100101000X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000000010000000  0X1101000X1XXXX01");
    apply_vector ( 24'b111001011000000010000000,17'b0X1101000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100000010000010  110011000X0XXXX00");
    apply_vector ( 24'b010001010100000010000010,17'b110011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100000010000000  0X1011000X0XXXX00");
    apply_vector ( 24'b111001011100000010000000,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010000010000001  100111000X0XXXX00");
    apply_vector ( 24'b001001010010000010000001,17'b100111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111001011010000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110000010000001  110000100X0XXXX00");
    apply_vector ( 24'b010001010110000010000001,17'b110000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110000010000000  0X1000100X0XXXX00");
    apply_vector ( 24'b111001011110000010000000,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001000010000000  100100100X0XXXX00");
    apply_vector ( 24'b001001010001000010000000,17'b100100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001000010000000  0X1100100X1000011");
    apply_vector ( 24'b111001011001000010000000,17'b0X1100100X1000011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101000010000011  110010100X0000010");
    apply_vector ( 24'b010001010101000010000011,17'b110010100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101000010000000  0X1010100X0000010");
    apply_vector ( 24'b111001011101000010000000,17'b0X1010100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011000010000001  100110100X0000010");
    apply_vector ( 24'b001001010011000010000001,17'b100110100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011000010000000  0X1110100X0000010");
    apply_vector ( 24'b111001011011000010000000,17'b0X1110100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111000010000001  110001100X0000010");
    apply_vector ( 24'b010001010111000010000001,17'b110001100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111000010000000  0X1001100X0000010");
    apply_vector ( 24'b111001011111000010000000,17'b0X1001100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000000010000000  101101000X0000010");
    apply_vector ( 24'b001011010000000010000000,17'b101101000X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000000010000000  0X0011000X1000010");
    apply_vector ( 24'b111011011000000010000000,17'b0X0011000X1000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100000010000010  111011000X0000010");
    apply_vector ( 24'b010011010100000010000010,17'b111011000X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100000010000001  0X0111000X0000010");
    apply_vector ( 24'b111011011100000010000001,17'b0X0111000X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010000010000001  101111000X0000010");
    apply_vector ( 24'b001011010010000010000001,17'b101111000X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010000010000000  0X0000100X0000010");
    apply_vector ( 24'b111011011010000010000000,17'b0X0000100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110000010000001  111000100X0000010");
    apply_vector ( 24'b010011010110000010000001,17'b111000100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110000010000000  0X0100100X0000010");
    apply_vector ( 24'b111011011110000010000000,17'b0X0100100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001000010000000  101100100X0000010");
    apply_vector ( 24'b001011010001000010000000,17'b101100100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001000010000000  0X0010100X1XXXX01");
    apply_vector ( 24'b111011011001000010000000,17'b0X0010100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101000010000011  111010100X0XXXX00");
    apply_vector ( 24'b010011010101000010000011,17'b111010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101000010000001  0X0110100X0XXXX00");
    apply_vector ( 24'b111011011101000010000001,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011000010000001  101110100X0XXXX00");
    apply_vector ( 24'b001011010011000010000001,17'b101110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011000010000000  0X0001100X0XXXX00");
    apply_vector ( 24'b111011011011000010000000,17'b0X0001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111000010000001  111001100X0XXXX00");
    apply_vector ( 24'b010011010111000010000001,17'b111001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111000010000000  0X0101100X0XXXX00");
    apply_vector ( 24'b111011011111000010000000,17'b0X0101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000000010000000  100011000X0XXXX00");
    apply_vector ( 24'b001000110000000010000000,17'b100011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000000010000000  0X1011000X1000011");
    apply_vector ( 24'b111000111000000010000000,17'b0X1011000X1000011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100000010000010  110111000X0000010");
    apply_vector ( 24'b010000110100000010000010,17'b110111000X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100000010000000  0X1111000X0000010");
    apply_vector ( 24'b111000111100000010000000,17'b0X1111000X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010000010000000  100000100X0000010");
    apply_vector ( 24'b001000110010000010000000,17'b100000100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010000010000001  0X1000100X0000010");
    apply_vector ( 24'b111000111010000010000001,17'b0X1000100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110000010000001  110100100X0000010");
    apply_vector ( 24'b010000110110000010000001,17'b110100100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110000010000000  0X1100100X0000010");
    apply_vector ( 24'b111000111110000010000000,17'b0X1100100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001000010000000  100010100X0000010");
    apply_vector ( 24'b001000110001000010000000,17'b100010100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001000010000000  0X1010100X1011011");
    apply_vector ( 24'b111000111001000010000000,17'b0X1010100X1011011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101000010000011  110110100X0011010");
    apply_vector ( 24'b010000110101000010000011,17'b110110100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101000010000000  0X1110100X0011010");
    apply_vector ( 24'b111000111101000010000000,17'b0X1110100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011000010000000  100001100X0011010");
    apply_vector ( 24'b001000110011000010000000,17'b100001100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011000010000001  0X1001100X0011010");
    apply_vector ( 24'b111000111011000010000001,17'b0X1001100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111000010000001  110101100X0011010");
    apply_vector ( 24'b010000110111000010000001,17'b110101100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111000010000000  0X1101100X0011010");
    apply_vector ( 24'b111000111111000010000000,17'b0X1101100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000000010000000  101011000X0011010");
    apply_vector ( 24'b001010110000000010000000,17'b101011000X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000000010000000  0X0111000X1XXXX01");
    apply_vector ( 24'b111010111000000010000000,17'b0X0111000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100000010000010  111111000X0XXXX00");
    apply_vector ( 24'b010010110100000010000010,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100000010000001  0X0000100X0XXXX00");
    apply_vector ( 24'b111010111100000010000001,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010000010000000  101000100X0XXXX00");
    apply_vector ( 24'b001010110010000010000000,17'b101000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010000010000001  0X0100100X0XXXX00");
    apply_vector ( 24'b111010111010000010000001,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110000010000001  111100100X0XXXX00");
    apply_vector ( 24'b010010110110000010000001,17'b111100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110000010000000  0X0010100X0XXXX00");
    apply_vector ( 24'b111010111110000010000000,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001000010000000  101010100X0XXXX00");
    apply_vector ( 24'b001010110001000010000000,17'b101010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001000010000000  0X0110100X1XXXX01");
    apply_vector ( 24'b111010111001000010000000,17'b0X0110100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101000010000011  111110100X0XXXX00");
    apply_vector ( 24'b010010110101000010000011,17'b111110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101000010000001  0X0001100X0XXXX00");
    apply_vector ( 24'b111010111101000010000001,17'b0X0001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011000010000000  101001100X0XXXX00");
    apply_vector ( 24'b001010110011000010000000,17'b101001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011000010000001  0X0101100X0XXXX00");
    apply_vector ( 24'b111010111011000010000001,17'b0X0101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111000010000001  111101100X0XXXX00");
    apply_vector ( 24'b010010110111000010000001,17'b111101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111000010000000  0X0011100X0XXXX00");
    apply_vector ( 24'b111010111111000010000000,17'b0X0011100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000000010000000  100111000X0XXXX00");
    apply_vector ( 24'b001001110000000010000000,17'b100111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000000010000000  0X1111000X1110111");
    apply_vector ( 24'b111001111000000010000000,17'b0X1111000X1110111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100000010000010  110000100X0110110");
    apply_vector ( 24'b010001110100000010000010,17'b110000100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100000010000000  0X1000100X0110110");
    apply_vector ( 24'b111001111100000010000000,17'b0X1000100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010000010000001  100100100X0110110");
    apply_vector ( 24'b001001110010000010000001,17'b100100100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010000010000001  0X1100100X0110110");
    apply_vector ( 24'b111001111010000010000001,17'b0X1100100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110000010000001  110010100X0110110");
    apply_vector ( 24'b010001110110000010000001,17'b110010100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110000010000000  0X1010100X0110110");
    apply_vector ( 24'b111001111110000010000000,17'b0X1010100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001000010000000  100110100X0110110");
    apply_vector ( 24'b001001110001000010000000,17'b100110100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001000010000000  0X1110100X1XXXX01");
    apply_vector ( 24'b111001111001000010000000,17'b0X1110100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101000010000011  110001100X0XXXX00");
    apply_vector ( 24'b010001110101000010000011,17'b110001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101000010000000  0X1001100X0XXXX00");
    apply_vector ( 24'b111001111101000010000000,17'b0X1001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011000010000001  100101100X0XXXX00");
    apply_vector ( 24'b001001110011000010000001,17'b100101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011000010000001  0X1101100X0XXXX00");
    apply_vector ( 24'b111001111011000010000001,17'b0X1101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111000010000001  110011100X0XXXX00");
    apply_vector ( 24'b010001110111000010000001,17'b110011100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111000010000000  0X1011100X0XXXX00");
    apply_vector ( 24'b111001111111000010000000,17'b0X1011100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000000010000000  101111000X0XXXX00");
    apply_vector ( 24'b001011110000000010000000,17'b101111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000000010000000  0X0000100X1000011");
    apply_vector ( 24'b111011111000000010000000,17'b0X0000100X1000011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100000010000010  111000100X0000010");
    apply_vector ( 24'b010011110100000010000010,17'b111000100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100000010000001  0X0100100X0000010");
    apply_vector ( 24'b111011111100000010000001,17'b0X0100100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010000010000001  101100100X0000010");
    apply_vector ( 24'b001011110010000010000001,17'b101100100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010000010000001  0X0010100X0000010");
    apply_vector ( 24'b111011111010000010000001,17'b0X0010100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110000010000001  111010100X0000010");
    apply_vector ( 24'b010011110110000010000001,17'b111010100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110000010000000  0X0110100X0000010");
    apply_vector ( 24'b111011111110000010000000,17'b0X0110100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001000010000000  101110100X0000010");
    apply_vector ( 24'b001011110001000010000000,17'b101110100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001000010000000  0X0001100X1110011");
    apply_vector ( 24'b111011111001000010000000,17'b0X0001100X1110011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101000010000011  111001100X0110010");
    apply_vector ( 24'b010011110101000010000011,17'b111001100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101000010000001  0X0101100X0110010");
    apply_vector ( 24'b111011111101000010000001,17'b0X0101100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011000010000001  101101100X0110010");
    apply_vector ( 24'b001011110011000010000001,17'b101101100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011000010000001  0X0011100X0110010");
    apply_vector ( 24'b111011111011000010000001,17'b0X0011100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111000010000001  111011100X0110010");
    apply_vector ( 24'b010011110111000010000001,17'b111011100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111000010000000  0X0111100X0110010");
    apply_vector ( 24'b111011111111000010000000,17'b0X0111100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100000000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000000010000000  101000000X0110010");
    apply_vector ( 24'b001100000000000010000000,17'b101000000X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000000010000000  0X0100000X1XXXX01");
    apply_vector ( 24'b111100001000000010000000,17'b0X0100000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100000010000010  111100000X0XXXX00");
    apply_vector ( 24'b010100000100000010000010,17'b111100000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100000010000000  0X0010000X0XXXX00");
    apply_vector ( 24'b111100001100000010000000,17'b0X0010000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010000010000000  101010000X0XXXX00");
    apply_vector ( 24'b001100000010000010000000,17'b101010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010000010000000  0X0110000X0XXXX00");
    apply_vector ( 24'b111100001010000010000000,17'b0X0110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110000010000000  111110000X0XXXX00");
    apply_vector ( 24'b010100000110000010000000,17'b111110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110000010000001  0X0001000X0XXXX00");
    apply_vector ( 24'b111100001110000010000001,17'b0X0001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001000010000000  101001000X0XXXX00");
    apply_vector ( 24'b001100000001000010000000,17'b101001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001000010000000  0X0101000X1XXXX01");
    apply_vector ( 24'b111100001001000010000000,17'b0X0101000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101000010000011  111101000X0XXXX00");
    apply_vector ( 24'b010100000101000010000011,17'b111101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101000010000000  0X0011000X0XXXX00");
    apply_vector ( 24'b111100001101000010000000,17'b0X0011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011000010000000  101011000X0XXXX00");
    apply_vector ( 24'b001100000011000010000000,17'b101011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011000010000000  0X0111000X0XXXX00");
    apply_vector ( 24'b111100001011000010000000,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111000010000000  111111000X0XXXX00");
    apply_vector ( 24'b010100000111000010000000,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111000010000001  0X0000100X0XXXX00");
    apply_vector ( 24'b111100001111000010000001,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110000000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000000010000000  100100000X0XXXX00");
    apply_vector ( 24'b001110000000000010000000,17'b100100000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110001000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000000010000000  0X1100000X1001111");
    apply_vector ( 24'b111110001000000010000000,17'b0X1100000X1001111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100000010000010  110010000X0001110");
    apply_vector ( 24'b010110000100000010000010,17'b110010000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100000010000001  0X1010000X0001110");
    apply_vector ( 24'b111110001100000010000001,17'b0X1010000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010000010000000  100110000X0001110");
    apply_vector ( 24'b001110000010000010000000,17'b100110000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010000010000000  0X1110000X0001110");
    apply_vector ( 24'b111110001010000010000000,17'b0X1110000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110000010000000  110001000X0001110");
    apply_vector ( 24'b010110000110000010000000,17'b110001000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110000010000001  0X1001000X0001110");
    apply_vector ( 24'b111110001110000010000001,17'b0X1001000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001000010000000  100101000X0001110");
    apply_vector ( 24'b001110000001000010000000,17'b100101000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001000010000000  0X1101000X1100011");
    apply_vector ( 24'b111110001001000010000000,17'b0X1101000X1100011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101000010000011  110011000X0100010");
    apply_vector ( 24'b010110000101000010000011,17'b110011000X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101000010000001  0X1011000X0100010");
    apply_vector ( 24'b111110001101000010000001,17'b0X1011000X0100010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011000010000000  100111000X0100010");
    apply_vector ( 24'b001110000011000010000000,17'b100111000X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011000010000000  0X1111000X0100010");
    apply_vector ( 24'b111110001011000010000000,17'b0X1111000X0100010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111000010000000  110000100X0100010");
    apply_vector ( 24'b010110000111000010000000,17'b110000100X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111000010000001  0X1000100X0100010");
    apply_vector ( 24'b111110001111000010000001,17'b0X1000100X0100010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101000000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000000010000000  101100000X0100010");
    apply_vector ( 24'b001101000000000010000000,17'b101100000X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000000010000000  0X0010000X1XXXX01");
    apply_vector ( 24'b111101001000000010000000,17'b0X0010000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100000010000010  111010000X0XXXX00");
    apply_vector ( 24'b010101000100000010000010,17'b111010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100000010000000  0X0110000X0XXXX00");
    apply_vector ( 24'b111101001100000010000000,17'b0X0110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010000010000001  101110000X0XXXX00");
    apply_vector ( 24'b001101000010000010000001,17'b101110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010000010000000  0X0001000X0XXXX00");
    apply_vector ( 24'b111101001010000010000000,17'b0X0001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110000010000000  111001000X0XXXX00");
    apply_vector ( 24'b010101000110000010000000,17'b111001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110000010000001  0X0101000X0XXXX00");
    apply_vector ( 24'b111101001110000010000001,17'b0X0101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001000010000000  101101000X0XXXX00");
    apply_vector ( 24'b001101000001000010000000,17'b101101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001000010000000  0X0011000X1001011");
    apply_vector ( 24'b111101001001000010000000,17'b0X0011000X1001011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101000010000011  111011000X0001010");
    apply_vector ( 24'b010101000101000010000011,17'b111011000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101000010000000  0X0111000X0001010");
    apply_vector ( 24'b111101001101000010000000,17'b0X0111000X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011000010000001  101111000X0001010");
    apply_vector ( 24'b001101000011000010000001,17'b101111000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011000010000000  0X0000100X0001010");
    apply_vector ( 24'b111101001011000010000000,17'b0X0000100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111000010000000  111000100X0001010");
    apply_vector ( 24'b010101000111000010000000,17'b111000100X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111000010000001  0X0100100X0001010");
    apply_vector ( 24'b111101001111000010000001,17'b0X0100100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111000000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000000010000000  100010000X0001010");
    apply_vector ( 24'b001111000000000010000000,17'b100010000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000000010000000  0X1010000X1XXXX01");
    apply_vector ( 24'b111111001000000010000000,17'b0X1010000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100000010000010  110110000X0XXXX00");
    apply_vector ( 24'b010111000100000010000010,17'b110110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100000010000001  0X1110000X0XXXX00");
    apply_vector ( 24'b111111001100000010000001,17'b0X1110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010000010000001  100001000X0XXXX00");
    apply_vector ( 24'b001111000010000010000001,17'b100001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010000010000000  0X1001000X0XXXX00");
    apply_vector ( 24'b111111001010000010000000,17'b0X1001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110000010000000  110101000X0XXXX00");
    apply_vector ( 24'b010111000110000010000000,17'b110101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110000010000001  0X1101000X0XXXX00");
    apply_vector ( 24'b111111001110000010000001,17'b0X1101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001000010000000  100011000X0XXXX00");
    apply_vector ( 24'b001111000001000010000000,17'b100011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001000010000000  0X1011000X1XXXX01");
    apply_vector ( 24'b111111001001000010000000,17'b0X1011000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101000010000011  110111000X0XXXX00");
    apply_vector ( 24'b010111000101000010000011,17'b110111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101000010000001  0X1111000X0XXXX00");
    apply_vector ( 24'b111111001101000010000001,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011000010000001  100000100X0XXXX00");
    apply_vector ( 24'b001111000011000010000001,17'b100000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011000010000000  0X1000100X0XXXX00");
    apply_vector ( 24'b111111001011000010000000,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111000010000000  110100100X0XXXX00");
    apply_vector ( 24'b010111000111000010000000,17'b110100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111000010000001  0X1100100X0XXXX00");
    apply_vector ( 24'b111111001111000010000001,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100100000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000000010000000  101010000X0XXXX00");
    apply_vector ( 24'b001100100000000010000000,17'b101010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000000010000000  0X0110000X1111011");
    apply_vector ( 24'b111100101000000010000000,17'b0X0110000X1111011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100000010000010  111110000X0111010");
    apply_vector ( 24'b010100100100000010000010,17'b111110000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100000010000000  0X0001000X0111010");
    apply_vector ( 24'b111100101100000010000000,17'b0X0001000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010000010000000  101001000X0111010");
    apply_vector ( 24'b001100100010000010000000,17'b101001000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010000010000001  0X0101000X0111010");
    apply_vector ( 24'b111100101010000010000001,17'b0X0101000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110000010000000  111101000X0111010");
    apply_vector ( 24'b010100100110000010000000,17'b111101000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110000010000001  0X0011000X0111010");
    apply_vector ( 24'b111100101110000010000001,17'b0X0011000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100100001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001000010000000  101011000X0111010");
    apply_vector ( 24'b001100100001000010000000,17'b101011000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001000010000000  0X0111000X1011011");
    apply_vector ( 24'b111100101001000010000000,17'b0X0111000X1011011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101000010000011  111111000X0011010");
    apply_vector ( 24'b010100100101000010000011,17'b111111000X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101000010000000  0X0000100X0011010");
    apply_vector ( 24'b111100101101000010000000,17'b0X0000100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011000010000000  101000100X0011010");
    apply_vector ( 24'b001100100011000010000000,17'b101000100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011000010000001  0X0100100X0011010");
    apply_vector ( 24'b111100101011000010000001,17'b0X0100100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111000010000000  111100100X0011010");
    apply_vector ( 24'b010100100111000010000000,17'b111100100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111000010000001  0X0010100X0011010");
    apply_vector ( 24'b111100101111000010000001,17'b0X0010100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110100000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000000010000000  100110000X0011010");
    apply_vector ( 24'b001110100000000010000000,17'b100110000X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000000010000000  0X1110000X1XXXX01");
    apply_vector ( 24'b111110101000000010000000,17'b0X1110000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100000010000010  110001000X0XXXX00");
    apply_vector ( 24'b010110100100000010000010,17'b110001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100000010000001  0X1001000X0XXXX00");
    apply_vector ( 24'b111110101100000010000001,17'b0X1001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010000010000000  100101000X0XXXX00");
    apply_vector ( 24'b001110100010000010000000,17'b100101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010000010000001  0X1101000X0XXXX00");
    apply_vector ( 24'b111110101010000010000001,17'b0X1101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110000010000000  110011000X0XXXX00");
    apply_vector ( 24'b010110100110000010000000,17'b110011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110000010000001  0X1011000X0XXXX00");
    apply_vector ( 24'b111110101110000010000001,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110100001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001000010000000  100111000X0XXXX00");
    apply_vector ( 24'b001110100001000010000000,17'b100111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110101001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001000010000000  0X1111000X1XXXX01");
    apply_vector ( 24'b111110101001000010000000,17'b0X1111000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101000010000011  110000100X0XXXX00");
    apply_vector ( 24'b010110100101000010000011,17'b110000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101000010000001  0X1000100X0XXXX00");
    apply_vector ( 24'b111110101101000010000001,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011000010000000  100100100X0XXXX00");
    apply_vector ( 24'b001110100011000010000000,17'b100100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011000010000001  0X1100100X0XXXX00");
    apply_vector ( 24'b111110101011000010000001,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111000010000000  110010100X0XXXX00");
    apply_vector ( 24'b010110100111000010000000,17'b110010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111000010000001  0X1010100X0XXXX00");
    apply_vector ( 24'b111110101111000010000001,17'b0X1010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101100000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000000010000000  101110000X0XXXX00");
    apply_vector ( 24'b001101100000000010000000,17'b101110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000000010000000  0X0001000X1111011");
    apply_vector ( 24'b111101101000000010000000,17'b0X0001000X1111011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100000010000010  111001000X0111010");
    apply_vector ( 24'b010101100100000010000010,17'b111001000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100000010000000  0X0101000X0111010");
    apply_vector ( 24'b111101101100000010000000,17'b0X0101000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010000010000001  101101000X0111010");
    apply_vector ( 24'b001101100010000010000001,17'b101101000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010000010000001  0X0011000X0111010");
    apply_vector ( 24'b111101101010000010000001,17'b0X0011000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110000010000000  111011000X0111010");
    apply_vector ( 24'b010101100110000010000000,17'b111011000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110000010000001  0X0111000X0111010");
    apply_vector ( 24'b111101101110000010000001,17'b0X0111000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101100001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001000010000000  101111000X0111010");
    apply_vector ( 24'b001101100001000010000000,17'b101111000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001000010000000  0X0000100X1XXXX01");
    apply_vector ( 24'b111101101001000010000000,17'b0X0000100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101000010000011  111000100X0XXXX00");
    apply_vector ( 24'b010101100101000010000011,17'b111000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101000010000000  0X0100100X0XXXX00");
    apply_vector ( 24'b111101101101000010000000,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011000010000001  101100100X0XXXX00");
    apply_vector ( 24'b001101100011000010000001,17'b101100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011000010000001  0X0010100X0XXXX00");
    apply_vector ( 24'b111101101011000010000001,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111000010000000  111010100X0XXXX00");
    apply_vector ( 24'b010101100111000010000000,17'b111010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111000010000001  0X0110100X0XXXX00");
    apply_vector ( 24'b111101101111000010000001,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111100000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000000010000000  100001000X0XXXX00");
    apply_vector ( 24'b001111100000000010000000,17'b100001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000000010000000  0X1001000X1111011");
    apply_vector ( 24'b111111101000000010000000,17'b0X1001000X1111011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100000010000010  110101000X0111010");
    apply_vector ( 24'b010111100100000010000010,17'b110101000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100000010000001  0X1101000X0111010");
    apply_vector ( 24'b111111101100000010000001,17'b0X1101000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010000010000001  100011000X0111010");
    apply_vector ( 24'b001111100010000010000001,17'b100011000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010000010000001  0X1011000X0111010");
    apply_vector ( 24'b111111101010000010000001,17'b0X1011000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110000010000000  110111000X0111010");
    apply_vector ( 24'b010111100110000010000000,17'b110111000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110000010000001  0X1111000X0111010");
    apply_vector ( 24'b111111101110000010000001,17'b0X1111000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111100001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001000010000000  100000100X0111010");
    apply_vector ( 24'b001111100001000010000000,17'b100000100X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001000010000000  0X1000100X1111011");
    apply_vector ( 24'b111111101001000010000000,17'b0X1000100X1111011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101000010000011  110100100X0111010");
    apply_vector ( 24'b010111100101000010000011,17'b110100100X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101000010000001  0X1100100X0111010");
    apply_vector ( 24'b111111101101000010000001,17'b0X1100100X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011000010000001  100010100X0111010");
    apply_vector ( 24'b001111100011000010000001,17'b100010100X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011000010000001  0X1010100X0111010");
    apply_vector ( 24'b111111101011000010000001,17'b0X1010100X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111000010000000  110110100X0111010");
    apply_vector ( 24'b010111100111000010000000,17'b110110100X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111000010000001  0X1110100X0111010");
    apply_vector ( 24'b111111101111000010000001,17'b0X1110100X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000000010000000  101001000X0111010");
    apply_vector ( 24'b001100010000000010000000,17'b101001000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000000010000000  0X0101000X1111010");
    apply_vector ( 24'b111100011000000010000000,17'b0X0101000X1111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100000010000010  111101000X0111010");
    apply_vector ( 24'b010100010100000010000010,17'b111101000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100000010000000  0X0011000X0111010");
    apply_vector ( 24'b111100011100000010000000,17'b0X0011000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010000010000000  101011000X0111010");
    apply_vector ( 24'b001100010010000010000000,17'b101011000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010000010000000  0X0111000X0111010");
    apply_vector ( 24'b111100011010000010000000,17'b0X0111000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110000010000001  111111000X0111010");
    apply_vector ( 24'b010100010110000010000001,17'b111111000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110000010000001  0X0000100X0111010");
    apply_vector ( 24'b111100011110000010000001,17'b0X0000100X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001000010000000  101000100X0111010");
    apply_vector ( 24'b001100010001000010000000,17'b101000100X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001000010000000  0X0100100X1011011");
    apply_vector ( 24'b111100011001000010000000,17'b0X0100100X1011011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101000010000011  111100100X0011010");
    apply_vector ( 24'b010100010101000010000011,17'b111100100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101000010000000  0X0010100X0011010");
    apply_vector ( 24'b111100011101000010000000,17'b0X0010100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011000010000000  101010100X0011010");
    apply_vector ( 24'b001100010011000010000000,17'b101010100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011000010000000  0X0110100X0011010");
    apply_vector ( 24'b111100011011000010000000,17'b0X0110100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111000010000001  111110100X0011010");
    apply_vector ( 24'b010100010111000010000001,17'b111110100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111000010000001  0X0001100X0011010");
    apply_vector ( 24'b111100011111000010000001,17'b0X0001100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000000010000000  100101000X0011010");
    apply_vector ( 24'b001110010000000010000000,17'b100101000X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000000010000000  0X1101000X1XXXX01");
    apply_vector ( 24'b111110011000000010000000,17'b0X1101000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100000010000010  110011000X0XXXX00");
    apply_vector ( 24'b010110010100000010000010,17'b110011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100000010000001  0X1011000X0XXXX00");
    apply_vector ( 24'b111110011100000010000001,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010000010000000  100111000X0XXXX00");
    apply_vector ( 24'b001110010010000010000000,17'b100111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111110011010000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110000010000001  110000100X0XXXX00");
    apply_vector ( 24'b010110010110000010000001,17'b110000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110000010000001  0X1000100X0XXXX00");
    apply_vector ( 24'b111110011110000010000001,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001000010000000  100100100X0XXXX00");
    apply_vector ( 24'b001110010001000010000000,17'b100100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001000010000000  0X1100100X1XXXX01");
    apply_vector ( 24'b111110011001000010000000,17'b0X1100100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101000010000011  110010100X0XXXX00");
    apply_vector ( 24'b010110010101000010000011,17'b110010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101000010000001  0X1010100X0XXXX00");
    apply_vector ( 24'b111110011101000010000001,17'b0X1010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011000010000000  100110100X0XXXX00");
    apply_vector ( 24'b001110010011000010000000,17'b100110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011000010000000  0X1110100X0XXXX00");
    apply_vector ( 24'b111110011011000010000000,17'b0X1110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111000010000001  110001100X0XXXX00");
    apply_vector ( 24'b010110010111000010000001,17'b110001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111000010000001  0X1001100X0XXXX00");
    apply_vector ( 24'b111110011111000010000001,17'b0X1001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000000010000000  101101000X0XXXX00");
    apply_vector ( 24'b001101010000000010000000,17'b101101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000000010000000  0X0011000X1101011");
    apply_vector ( 24'b111101011000000010000000,17'b0X0011000X1101011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100000010000010  111011000X0101010");
    apply_vector ( 24'b010101010100000010000010,17'b111011000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100000010000000  0X0111000X0101010");
    apply_vector ( 24'b111101011100000010000000,17'b0X0111000X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010000010000001  101111000X0101010");
    apply_vector ( 24'b001101010010000010000001,17'b101111000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010000010000000  0X0000100X0101010");
    apply_vector ( 24'b111101011010000010000000,17'b0X0000100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110000010000001  111000100X0101010");
    apply_vector ( 24'b010101010110000010000001,17'b111000100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110000010000001  0X0100100X0101010");
    apply_vector ( 24'b111101011110000010000001,17'b0X0100100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001000010000000  101100100X0101010");
    apply_vector ( 24'b001101010001000010000000,17'b101100100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001000010000000  0X0010100X1XXXX01");
    apply_vector ( 24'b111101011001000010000000,17'b0X0010100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101000010000011  111010100X0XXXX00");
    apply_vector ( 24'b010101010101000010000011,17'b111010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101000010000000  0X0110100X0XXXX00");
    apply_vector ( 24'b111101011101000010000000,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011000010000001  101110100X0XXXX00");
    apply_vector ( 24'b001101010011000010000001,17'b101110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011000010000000  0X0001100X0XXXX00");
    apply_vector ( 24'b111101011011000010000000,17'b0X0001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111000010000001  111001100X0XXXX00");
    apply_vector ( 24'b010101010111000010000001,17'b111001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111000010000001  0X0101100X0XXXX00");
    apply_vector ( 24'b111101011111000010000001,17'b0X0101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000000010000000  100011000X0XXXX00");
    apply_vector ( 24'b001111010000000010000000,17'b100011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000000010000000  0X1011000X1000011");
    apply_vector ( 24'b111111011000000010000000,17'b0X1011000X1000011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100000010000010  110111000X0000010");
    apply_vector ( 24'b010111010100000010000010,17'b110111000X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100000010000001  0X1111000X0000010");
    apply_vector ( 24'b111111011100000010000001,17'b0X1111000X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010000010000001  100000100X0000010");
    apply_vector ( 24'b001111010010000010000001,17'b100000100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010000010000000  0X1000100X0000010");
    apply_vector ( 24'b111111011010000010000000,17'b0X1000100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110000010000001  110100100X0000010");
    apply_vector ( 24'b010111010110000010000001,17'b110100100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110000010000001  0X1100100X0000010");
    apply_vector ( 24'b111111011110000010000001,17'b0X1100100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001000010000000  100010100X0000010");
    apply_vector ( 24'b001111010001000010000000,17'b100010100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001000010000000  0X1010100X1101111");
    apply_vector ( 24'b111111011001000010000000,17'b0X1010100X1101111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101000010000011  110110100X0101110");
    apply_vector ( 24'b010111010101000010000011,17'b110110100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101000010000001  0X1110100X0101110");
    apply_vector ( 24'b111111011101000010000001,17'b0X1110100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011000010000001  100001100X0101110");
    apply_vector ( 24'b001111010011000010000001,17'b100001100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011000010000000  0X1001100X0101110");
    apply_vector ( 24'b111111011011000010000000,17'b0X1001100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111000010000001  110101100X0101110");
    apply_vector ( 24'b010111010111000010000001,17'b110101100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111000010000001  0X1101100X0101110");
    apply_vector ( 24'b111111011111000010000001,17'b0X1101100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000000010000000  101011000X0101110");
    apply_vector ( 24'b001100110000000010000000,17'b101011000X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000000010000000  0X0111000X1XXXX01");
    apply_vector ( 24'b111100111000000010000000,17'b0X0111000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100000010000010  111111000X0XXXX00");
    apply_vector ( 24'b010100110100000010000010,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100000010000000  0X0000100X0XXXX00");
    apply_vector ( 24'b111100111100000010000000,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010000010000000  101000100X0XXXX00");
    apply_vector ( 24'b001100110010000010000000,17'b101000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010000010000001  0X0100100X0XXXX00");
    apply_vector ( 24'b111100111010000010000001,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110000010000001  111100100X0XXXX00");
    apply_vector ( 24'b010100110110000010000001,17'b111100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110000010000001  0X0010100X0XXXX00");
    apply_vector ( 24'b111100111110000010000001,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001000010000000  101010100X0XXXX00");
    apply_vector ( 24'b001100110001000010000000,17'b101010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001000010000000  0X0110100X1011010");
    apply_vector ( 24'b111100111001000010000000,17'b0X0110100X1011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101000010000011  111110100X0011010");
    apply_vector ( 24'b010100110101000010000011,17'b111110100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101000010000000  0X0001100X0011010");
    apply_vector ( 24'b111100111101000010000000,17'b0X0001100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011000010000000  101001100X0011010");
    apply_vector ( 24'b001100110011000010000000,17'b101001100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011000010000001  0X0101100X0011010");
    apply_vector ( 24'b111100111011000010000001,17'b0X0101100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111000010000001  111101100X0011010");
    apply_vector ( 24'b010100110111000010000001,17'b111101100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111000010000001  0X0011100X0011010");
    apply_vector ( 24'b111100111111000010000001,17'b0X0011100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000000010000000  100111000X0011010");
    apply_vector ( 24'b001110110000000010000000,17'b100111000X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000000010000000  0X1111000X1011011");
    apply_vector ( 24'b111110111000000010000000,17'b0X1111000X1011011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100000010000010  110000100X0011010");
    apply_vector ( 24'b010110110100000010000010,17'b110000100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100000010000001  0X1000100X0011010");
    apply_vector ( 24'b111110111100000010000001,17'b0X1000100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010000010000000  100100100X0011010");
    apply_vector ( 24'b001110110010000010000000,17'b100100100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010000010000001  0X1100100X0011010");
    apply_vector ( 24'b111110111010000010000001,17'b0X1100100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110000010000001  110010100X0011010");
    apply_vector ( 24'b010110110110000010000001,17'b110010100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110000010000001  0X1010100X0011010");
    apply_vector ( 24'b111110111110000010000001,17'b0X1010100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001000010000000  100110100X0011010");
    apply_vector ( 24'b001110110001000010000000,17'b100110100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001000010000000  0X1110100X1011011");
    apply_vector ( 24'b111110111001000010000000,17'b0X1110100X1011011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101000010000011  110001100X0011010");
    apply_vector ( 24'b010110110101000010000011,17'b110001100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101000010000001  0X1001100X0011010");
    apply_vector ( 24'b111110111101000010000001,17'b0X1001100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011000010000000  100101100X0011010");
    apply_vector ( 24'b001110110011000010000000,17'b100101100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011000010000001  0X1101100X0011010");
    apply_vector ( 24'b111110111011000010000001,17'b0X1101100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111000010000001  110011100X0011010");
    apply_vector ( 24'b010110110111000010000001,17'b110011100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111000010000001  0X1011100X0011010");
    apply_vector ( 24'b111110111111000010000001,17'b0X1011100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000000010000000  101111000X0011010");
    apply_vector ( 24'b001101110000000010000000,17'b101111000X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000000010000000  0X0000100X1XXXX01");
    apply_vector ( 24'b111101111000000010000000,17'b0X0000100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100000010000010  111000100X0XXXX00");
    apply_vector ( 24'b010101110100000010000010,17'b111000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100000010000000  0X0100100X0XXXX00");
    apply_vector ( 24'b111101111100000010000000,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010000010000001  101100100X0XXXX00");
    apply_vector ( 24'b001101110010000010000001,17'b101100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010000010000001  0X0010100X0XXXX00");
    apply_vector ( 24'b111101111010000010000001,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110000010000001  111010100X0XXXX00");
    apply_vector ( 24'b010101110110000010000001,17'b111010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110000010000001  0X0110100X0XXXX00");
    apply_vector ( 24'b111101111110000010000001,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001000010000000  101110100X0XXXX00");
    apply_vector ( 24'b001101110001000010000000,17'b101110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001000010000000  0X0001100X1011011");
    apply_vector ( 24'b111101111001000010000000,17'b0X0001100X1011011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101000010000011  111001100X0011010");
    apply_vector ( 24'b010101110101000010000011,17'b111001100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101000010000000  0X0101100X0011010");
    apply_vector ( 24'b111101111101000010000000,17'b0X0101100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011000010000001  101101100X0011010");
    apply_vector ( 24'b001101110011000010000001,17'b101101100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011000010000001  0X0011100X0011010");
    apply_vector ( 24'b111101111011000010000001,17'b0X0011100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111000010000001  111011100X0011010");
    apply_vector ( 24'b010101110111000010000001,17'b111011100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111000010000001  0X0111100X0011010");
    apply_vector ( 24'b111101111111000010000001,17'b0X0111100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000000010000000  100000100X0011010");
    apply_vector ( 24'b001111110000000010000000,17'b100000100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000000010000000  0X1000100X1XXXX01");
    apply_vector ( 24'b111111111000000010000000,17'b0X1000100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100000010000010  110100100X0XXXX00");
    apply_vector ( 24'b010111110100000010000010,17'b110100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100000010000001  0X1100100X0XXXX00");
    apply_vector ( 24'b111111111100000010000001,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010000010000001  100010100X0XXXX00");
    apply_vector ( 24'b001111110010000010000001,17'b100010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010000010000001  0X1010100X0XXXX00");
    apply_vector ( 24'b111111111010000010000001,17'b0X1010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110000010000001  110110100X0XXXX00");
    apply_vector ( 24'b010111110110000010000001,17'b110110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110000010000001  0X1110100X0XXXX00");
    apply_vector ( 24'b111111111110000010000001,17'b0X1110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001000010000000  100001100X0XXXX00");
    apply_vector ( 24'b001111110001000010000000,17'b100001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001000010000000  0X1001100X1XXXX01");
    apply_vector ( 24'b111111111001000010000000,17'b0X1001100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101000010000011  110101100X0XXXX00");
    apply_vector ( 24'b010111110101000010000011,17'b110101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101000010000001  0X1101100X0XXXX00");
    apply_vector ( 24'b111111111101000010000001,17'b0X1101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011000010000001  100011100X0XXXX00");
    apply_vector ( 24'b001111110011000010000001,17'b100011100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011000010000001  0X1011100X0XXXX00");
    apply_vector ( 24'b111111111011000010000001,17'b0X1011100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111000010000001  110111100X0XXXX00");
    apply_vector ( 24'b010111110111000010000001,17'b110111100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111000010000001  0X1111100X0XXXX00");
    apply_vector ( 24'b111111111111000010000001,17'b0X1111100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000000000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000000010000000  100000000X0XXXX00");
    apply_vector ( 24'b001000000000000010000000,17'b100000000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000000010000000  0X1000000X1111011");
    apply_vector ( 24'b111000001000000010000000,17'b0X1000000X1111011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100000010000010  110100000X0111010");
    apply_vector ( 24'b010000000100000010000010,17'b110100000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100000010000000  0X1100000X0111010");
    apply_vector ( 24'b111000001100000010000000,17'b0X1100000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010000010000000  100010000X0111010");
    apply_vector ( 24'b001000000010000010000000,17'b100010000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010000010000000  0X1010000X0111010");
    apply_vector ( 24'b111000001010000010000000,17'b0X1010000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110000010000000  110110000X0111010");
    apply_vector ( 24'b010000000110000010000000,17'b110110000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110000010000000  0X1110000X0111010");
    apply_vector ( 24'b111000001110000010000000,17'b0X1110000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001000010000001  100001000X0111010");
    apply_vector ( 24'b001000000001000010000001,17'b100001000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001000010000000  0X1001000X1XXXX01");
    apply_vector ( 24'b111000001001000010000000,17'b0X1001000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101000010000011  110101000X0XXXX00");
    apply_vector ( 24'b010000000101000010000011,17'b110101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101000010000000  0X1101000X0XXXX00");
    apply_vector ( 24'b111000001101000010000000,17'b0X1101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011000010000000  100011000X0XXXX00");
    apply_vector ( 24'b001000000011000010000000,17'b100011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011000010000000  0X1011000X0XXXX00");
    apply_vector ( 24'b111000001011000010000000,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111000010000000  110111000X0XXXX00");
    apply_vector ( 24'b010000000111000010000000,17'b110111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111000001111000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000000010000001  101000000X0XXXX00");
    apply_vector ( 24'b001010000000000010000001,17'b101000000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010001000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000000010000000  0X0100000X1010011");
    apply_vector ( 24'b111010001000000010000000,17'b0X0100000X1010011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100000010000010  111100000X0010010");
    apply_vector ( 24'b010010000100000010000010,17'b111100000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100000010000001  0X0010000X0010010");
    apply_vector ( 24'b111010001100000010000001,17'b0X0010000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010000010000000  101010000X0010010");
    apply_vector ( 24'b001010000010000010000000,17'b101010000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010000010000000  0X0110000X0010010");
    apply_vector ( 24'b111010001010000010000000,17'b0X0110000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110000010000000  111110000X0010010");
    apply_vector ( 24'b010010000110000010000000,17'b111110000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110000010000000  0X0001000X0010010");
    apply_vector ( 24'b111010001110000010000000,17'b0X0001000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001000010000001  101001000X0010010");
    apply_vector ( 24'b001010000001000010000001,17'b101001000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001000010000000  0X0101000X1100011");
    apply_vector ( 24'b111010001001000010000000,17'b0X0101000X1100011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101000010000011  111101000X0100010");
    apply_vector ( 24'b010010000101000010000011,17'b111101000X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101000010000001  0X0011000X0100010");
    apply_vector ( 24'b111010001101000010000001,17'b0X0011000X0100010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011000010000000  101011000X0100010");
    apply_vector ( 24'b001010000011000010000000,17'b101011000X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011000010000000  0X0111000X0100010");
    apply_vector ( 24'b111010001011000010000000,17'b0X0111000X0100010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111000010000000  111111000X0100010");
    apply_vector ( 24'b010010000111000010000000,17'b111111000X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111000010000000  0X0000100X0100010");
    apply_vector ( 24'b111010001111000010000000,17'b0X0000100X0100010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000000010000001  100100000X0100010");
    apply_vector ( 24'b001001000000000010000001,17'b100100000X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001001000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000000010000000  0X1100000X1XXXX01");
    apply_vector ( 24'b111001001000000010000000,17'b0X1100000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100000010000010  110010000X0XXXX00");
    apply_vector ( 24'b010001000100000010000010,17'b110010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100000010000000  0X1010000X0XXXX00");
    apply_vector ( 24'b111001001100000010000000,17'b0X1010000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010000010000001  100110000X0XXXX00");
    apply_vector ( 24'b001001000010000010000001,17'b100110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010000010000000  0X1110000X0XXXX00");
    apply_vector ( 24'b111001001010000010000000,17'b0X1110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110000010000000  110001000X0XXXX00");
    apply_vector ( 24'b010001000110000010000000,17'b110001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110000010000000  0X1001000X0XXXX00");
    apply_vector ( 24'b111001001110000010000000,17'b0X1001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001000010000001  100101000X0XXXX00");
    apply_vector ( 24'b001001000001000010000001,17'b100101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001000010000000  0X1101000X1001011");
    apply_vector ( 24'b111001001001000010000000,17'b0X1101000X1001011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101000010000011  110011000X0001010");
    apply_vector ( 24'b010001000101000010000011,17'b110011000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101000010000000  0X1011000X0001010");
    apply_vector ( 24'b111001001101000010000000,17'b0X1011000X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011000010000001  100111000X0001010");
    apply_vector ( 24'b001001000011000010000001,17'b100111000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011000010000000  0X1111000X0001010");
    apply_vector ( 24'b111001001011000010000000,17'b0X1111000X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111000010000000  110000100X0001010");
    apply_vector ( 24'b010001000111000010000000,17'b110000100X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001001111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111000010000000  0X1000100X0001010");
    apply_vector ( 24'b111001001111000010000000,17'b0X1000100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000000010000001  101100000X0001010");
    apply_vector ( 24'b001011000000000010000001,17'b101100000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011001000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000000010000000  0X0010000X1XXXX01");
    apply_vector ( 24'b111011001000000010000000,17'b0X0010000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100000010000010  111010000X0XXXX00");
    apply_vector ( 24'b010011000100000010000010,17'b111010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100000010000001  0X0110000X0XXXX00");
    apply_vector ( 24'b111011001100000010000001,17'b0X0110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010000010000001  101110000X0XXXX00");
    apply_vector ( 24'b001011000010000010000001,17'b101110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010000010000000  0X0001000X0XXXX00");
    apply_vector ( 24'b111011001010000010000000,17'b0X0001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110000010000000  111001000X0XXXX00");
    apply_vector ( 24'b010011000110000010000000,17'b111001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110000010000000  0X0101000X0XXXX00");
    apply_vector ( 24'b111011001110000010000000,17'b0X0101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001000010000001  101101000X0XXXX00");
    apply_vector ( 24'b001011000001000010000001,17'b101101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001000010000000  0X0011000X1XXXX01");
    apply_vector ( 24'b111011001001000010000000,17'b0X0011000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101000010000011  111011000X0XXXX00");
    apply_vector ( 24'b010011000101000010000011,17'b111011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101000010000001  0X0111000X0XXXX00");
    apply_vector ( 24'b111011001101000010000001,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011000010000001  101111000X0XXXX00");
    apply_vector ( 24'b001011000011000010000001,17'b101111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011000010000000  0X0000100X0XXXX00");
    apply_vector ( 24'b111011001011000010000000,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111000010000000  111000100X0XXXX00");
    apply_vector ( 24'b010011000111000010000000,17'b111000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111000010000000  0X0100100X0XXXX00");
    apply_vector ( 24'b111011001111000010000000,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000000010000001  100010000X0XXXX00");
    apply_vector ( 24'b001000100000000010000001,17'b100010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000101000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000000010000000  0X1010000X1100111");
    apply_vector ( 24'b111000101000000010000000,17'b0X1010000X1100111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100000010000010  110110000X0100110");
    apply_vector ( 24'b010000100100000010000010,17'b110110000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100000010000000  0X1110000X0100110");
    apply_vector ( 24'b111000101100000010000000,17'b0X1110000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010000010000000  100001000X0100110");
    apply_vector ( 24'b001000100010000010000000,17'b100001000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010000010000001  0X1001000X0100110");
    apply_vector ( 24'b111000101010000010000001,17'b0X1001000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110000010000000  110101000X0100110");
    apply_vector ( 24'b010000100110000010000000,17'b110101000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110000010000000  0X1101000X0100110");
    apply_vector ( 24'b111000101110000010000000,17'b0X1101000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001000010000001  100011000X0100110");
    apply_vector ( 24'b001000100001000010000001,17'b100011000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001000010000000  0X1011000X1010011");
    apply_vector ( 24'b111000101001000010000000,17'b0X1011000X1010011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101000010000011  110111000X0010010");
    apply_vector ( 24'b010000100101000010000011,17'b110111000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101000010000000  0X1111000X0010010");
    apply_vector ( 24'b111000101101000010000000,17'b0X1111000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011000010000000  100000100X0010010");
    apply_vector ( 24'b001000100011000010000000,17'b100000100X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011000010000001  0X1000100X0010010");
    apply_vector ( 24'b111000101011000010000001,17'b0X1000100X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111000010000000  110100100X0010010");
    apply_vector ( 24'b010000100111000010000000,17'b110100100X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111000010000000  0X1100100X0010010");
    apply_vector ( 24'b111000101111000010000000,17'b0X1100100X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000000010000001  101010000X0010010");
    apply_vector ( 24'b001010100000000010000001,17'b101010000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010101000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000000010000000  0X0110000X1010010");
    apply_vector ( 24'b111010101000000010000000,17'b0X0110000X1010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100000010000010  111110000X0010010");
    apply_vector ( 24'b010010100100000010000010,17'b111110000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100000010000001  0X0001000X0010010");
    apply_vector ( 24'b111010101100000010000001,17'b0X0001000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010000010000000  101001000X0010010");
    apply_vector ( 24'b001010100010000010000000,17'b101001000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010000010000001  0X0101000X0010010");
    apply_vector ( 24'b111010101010000010000001,17'b0X0101000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110000010000000  111101000X0010010");
    apply_vector ( 24'b010010100110000010000000,17'b111101000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010101110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110000010000000  0X0011000X0010010");
    apply_vector ( 24'b111010101110000010000000,17'b0X0011000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001000010000001  101011000X0010010");
    apply_vector ( 24'b001010100001000010000001,17'b101011000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010101001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001000010000000  0X0111000X1XXXX01");
    apply_vector ( 24'b111010101001000010000000,17'b0X0111000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101000010000011  111111000X0XXXX00");
    apply_vector ( 24'b010010100101000010000011,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101000010000001  0X0000100X0XXXX00");
    apply_vector ( 24'b111010101101000010000001,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011000010000000  101000100X0XXXX00");
    apply_vector ( 24'b001010100011000010000000,17'b101000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011000010000001  0X0100100X0XXXX00");
    apply_vector ( 24'b111010101011000010000001,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111000010000000  111100100X0XXXX00");
    apply_vector ( 24'b010010100111000010000000,17'b111100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010101111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111000010000000  0X0010100X0XXXX00");
    apply_vector ( 24'b111010101111000010000000,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000000010000001  100110000X0XXXX00");
    apply_vector ( 24'b001001100000000010000001,17'b100110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001101000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000000010000000  0X1110000X1010011");
    apply_vector ( 24'b111001101000000010000000,17'b0X1110000X1010011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100000010000010  110001000X0010010");
    apply_vector ( 24'b010001100100000010000010,17'b110001000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100000010000000  0X1001000X0010010");
    apply_vector ( 24'b111001101100000010000000,17'b0X1001000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010000010000001  100101000X0010010");
    apply_vector ( 24'b001001100010000010000001,17'b100101000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010000010000001  0X1101000X0010010");
    apply_vector ( 24'b111001101010000010000001,17'b0X1101000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110000010000000  110011000X0010010");
    apply_vector ( 24'b010001100110000010000000,17'b110011000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110000010000000  0X1011000X0010010");
    apply_vector ( 24'b111001101110000010000000,17'b0X1011000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001000010000001  100111000X0010010");
    apply_vector ( 24'b001001100001000010000001,17'b100111000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001000010000000  0X1111000X1XXXX01");
    apply_vector ( 24'b111001101001000010000000,17'b0X1111000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101000010000011  110000100X0XXXX00");
    apply_vector ( 24'b010001100101000010000011,17'b110000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101000010000000  0X1000100X0XXXX00");
    apply_vector ( 24'b111001101101000010000000,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011000010000001  100100100X0XXXX00");
    apply_vector ( 24'b001001100011000010000001,17'b100100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011000010000001  0X1100100X0XXXX00");
    apply_vector ( 24'b111001101011000010000001,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111000010000000  110010100X0XXXX00");
    apply_vector ( 24'b010001100111000010000000,17'b110010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001101111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111000010000000  0X1010100X0XXXX00");
    apply_vector ( 24'b111001101111000010000000,17'b0X1010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000000010000001  101110000X0XXXX00");
    apply_vector ( 24'b001011100000000010000001,17'b101110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011101000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000000010000000  0X0001000X1010011");
    apply_vector ( 24'b111011101000000010000000,17'b0X0001000X1010011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100000010000010  111001000X0010010");
    apply_vector ( 24'b010011100100000010000010,17'b111001000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100000010000001  0X0101000X0010010");
    apply_vector ( 24'b111011101100000010000001,17'b0X0101000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010000010000001  101101000X0010010");
    apply_vector ( 24'b001011100010000010000001,17'b101101000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010000010000001  0X0011000X0010010");
    apply_vector ( 24'b111011101010000010000001,17'b0X0011000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110000010000000  111011000X0010010");
    apply_vector ( 24'b010011100110000010000000,17'b111011000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110000010000000  0X0111000X0010010");
    apply_vector ( 24'b111011101110000010000000,17'b0X0111000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001000010000001  101111000X0010010");
    apply_vector ( 24'b001011100001000010000001,17'b101111000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001000010000000  0X0000100X1110011");
    apply_vector ( 24'b111011101001000010000000,17'b0X0000100X1110011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101000010000011  111000100X0110010");
    apply_vector ( 24'b010011100101000010000011,17'b111000100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101000010000001  0X0100100X0110010");
    apply_vector ( 24'b111011101101000010000001,17'b0X0100100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011000010000001  101100100X0110010");
    apply_vector ( 24'b001011100011000010000001,17'b101100100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011000010000001  0X0010100X0110010");
    apply_vector ( 24'b111011101011000010000001,17'b0X0010100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111000010000000  111010100X0110010");
    apply_vector ( 24'b010011100111000010000000,17'b111010100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111000010000000  0X0110100X0110010");
    apply_vector ( 24'b111011101111000010000000,17'b0X0110100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000000010000001  100001000X0110010");
    apply_vector ( 24'b001000010000000010000001,17'b100001000X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000000010000000  0X1001000X1XXXX01");
    apply_vector ( 24'b111000011000000010000000,17'b0X1001000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100000010000010  110101000X0XXXX00");
    apply_vector ( 24'b010000010100000010000010,17'b110101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100000010000000  0X1101000X0XXXX00");
    apply_vector ( 24'b111000011100000010000000,17'b0X1101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010000010000000  100011000X0XXXX00");
    apply_vector ( 24'b001000010010000010000000,17'b100011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010000010000000  0X1011000X0XXXX00");
    apply_vector ( 24'b111000011010000010000000,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110000010000001  110111000X0XXXX00");
    apply_vector ( 24'b010000010110000010000001,17'b110111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111000011110000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001000010000001  100000100X0XXXX00");
    apply_vector ( 24'b001000010001000010000001,17'b100000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001000010000000  0X1000100X1000111");
    apply_vector ( 24'b111000011001000010000000,17'b0X1000100X1000111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101000010000011  110100100X0000110");
    apply_vector ( 24'b010000010101000010000011,17'b110100100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101000010000000  0X1100100X0000110");
    apply_vector ( 24'b111000011101000010000000,17'b0X1100100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011000010000000  100010100X0000110");
    apply_vector ( 24'b001000010011000010000000,17'b100010100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011000010000000  0X1010100X0000110");
    apply_vector ( 24'b111000011011000010000000,17'b0X1010100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111000010000001  110110100X0000110");
    apply_vector ( 24'b010000010111000010000001,17'b110110100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111000010000000  0X1110100X0000110");
    apply_vector ( 24'b111000011111000010000000,17'b0X1110100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000000010000001  101001000X0000110");
    apply_vector ( 24'b001010010000000010000001,17'b101001000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000000010000000  0X0101000X1XXXX01");
    apply_vector ( 24'b111010011000000010000000,17'b0X0101000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100000010000010  111101000X0XXXX00");
    apply_vector ( 24'b010010010100000010000010,17'b111101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100000010000001  0X0011000X0XXXX00");
    apply_vector ( 24'b111010011100000010000001,17'b0X0011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010000010000000  101011000X0XXXX00");
    apply_vector ( 24'b001010010010000010000000,17'b101011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010000010000000  0X0111000X0XXXX00");
    apply_vector ( 24'b111010011010000010000000,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110000010000001  111111000X0XXXX00");
    apply_vector ( 24'b010010010110000010000001,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110000010000000  0X0000100X0XXXX00");
    apply_vector ( 24'b111010011110000010000000,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001000010000001  101000100X0XXXX00");
    apply_vector ( 24'b001010010001000010000001,17'b101000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001000010000000  0X0100100X1XXXX01");
    apply_vector ( 24'b111010011001000010000000,17'b0X0100100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101000010000011  111100100X0XXXX00");
    apply_vector ( 24'b010010010101000010000011,17'b111100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101000010000001  0X0010100X0XXXX00");
    apply_vector ( 24'b111010011101000010000001,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011000010000000  101010100X0XXXX00");
    apply_vector ( 24'b001010010011000010000000,17'b101010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011000010000000  0X0110100X0XXXX00");
    apply_vector ( 24'b111010011011000010000000,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111000010000001  111110100X0XXXX00");
    apply_vector ( 24'b010010010111000010000001,17'b111110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111000010000000  0X0001100X0XXXX00");
    apply_vector ( 24'b111010011111000010000000,17'b0X0001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000000010000001  100101000X0XXXX00");
    apply_vector ( 24'b001001010000000010000001,17'b100101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000000010000000  0X1101000X1101011");
    apply_vector ( 24'b111001011000000010000000,17'b0X1101000X1101011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100000010000010  110011000X0101010");
    apply_vector ( 24'b010001010100000010000010,17'b110011000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100000010000000  0X1011000X0101010");
    apply_vector ( 24'b111001011100000010000000,17'b0X1011000X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010000010000001  100111000X0101010");
    apply_vector ( 24'b001001010010000010000001,17'b100111000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010000010000000  0X1111000X0101010");
    apply_vector ( 24'b111001011010000010000000,17'b0X1111000X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110000010000001  110000100X0101010");
    apply_vector ( 24'b010001010110000010000001,17'b110000100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110000010000000  0X1000100X0101010");
    apply_vector ( 24'b111001011110000010000000,17'b0X1000100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001000010000001  100100100X0101010");
    apply_vector ( 24'b001001010001000010000001,17'b100100100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001000010000000  0X1100100X1XXXX01");
    apply_vector ( 24'b111001011001000010000000,17'b0X1100100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101000010000011  110010100X0XXXX00");
    apply_vector ( 24'b010001010101000010000011,17'b110010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101000010000000  0X1010100X0XXXX00");
    apply_vector ( 24'b111001011101000010000000,17'b0X1010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011000010000001  100110100X0XXXX00");
    apply_vector ( 24'b001001010011000010000001,17'b100110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011000010000000  0X1110100X0XXXX00");
    apply_vector ( 24'b111001011011000010000000,17'b0X1110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111000010000001  110001100X0XXXX00");
    apply_vector ( 24'b010001010111000010000001,17'b110001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111000010000000  0X1001100X0XXXX00");
    apply_vector ( 24'b111001011111000010000000,17'b0X1001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000000010000001  101101000X0XXXX00");
    apply_vector ( 24'b001011010000000010000001,17'b101101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000000010000000  0X0011000X1000011");
    apply_vector ( 24'b111011011000000010000000,17'b0X0011000X1000011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100000010000010  111011000X0000010");
    apply_vector ( 24'b010011010100000010000010,17'b111011000X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100000010000001  0X0111000X0000010");
    apply_vector ( 24'b111011011100000010000001,17'b0X0111000X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010000010000001  101111000X0000010");
    apply_vector ( 24'b001011010010000010000001,17'b101111000X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010000010000000  0X0000100X0000010");
    apply_vector ( 24'b111011011010000010000000,17'b0X0000100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110000010000001  111000100X0000010");
    apply_vector ( 24'b010011010110000010000001,17'b111000100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110000010000000  0X0100100X0000010");
    apply_vector ( 24'b111011011110000010000000,17'b0X0100100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001000010000001  101100100X0000010");
    apply_vector ( 24'b001011010001000010000001,17'b101100100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001000010000000  0X0010100X1110011");
    apply_vector ( 24'b111011011001000010000000,17'b0X0010100X1110011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101000010000011  111010100X0110010");
    apply_vector ( 24'b010011010101000010000011,17'b111010100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101000010000001  0X0110100X0110010");
    apply_vector ( 24'b111011011101000010000001,17'b0X0110100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011000010000001  101110100X0110010");
    apply_vector ( 24'b001011010011000010000001,17'b101110100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011000010000000  0X0001100X0110010");
    apply_vector ( 24'b111011011011000010000000,17'b0X0001100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111000010000001  111001100X0110010");
    apply_vector ( 24'b010011010111000010000001,17'b111001100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111000010000000  0X0101100X0110010");
    apply_vector ( 24'b111011011111000010000000,17'b0X0101100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000000010000001  100011000X0110010");
    apply_vector ( 24'b001000110000000010000001,17'b100011000X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000000010000000  0X1011000X1XXXX01");
    apply_vector ( 24'b111000111000000010000000,17'b0X1011000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100000010000010  110111000X0XXXX00");
    apply_vector ( 24'b010000110100000010000010,17'b110111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111000111100000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010000010000000  100000100X0XXXX00");
    apply_vector ( 24'b001000110010000010000000,17'b100000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010000010000001  0X1000100X0XXXX00");
    apply_vector ( 24'b111000111010000010000001,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110000010000001  110100100X0XXXX00");
    apply_vector ( 24'b010000110110000010000001,17'b110100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110000010000000  0X1100100X0XXXX00");
    apply_vector ( 24'b111000111110000010000000,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001000010000001  100010100X0XXXX00");
    apply_vector ( 24'b001000110001000010000001,17'b100010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001000010000000  0X1010100X1XXXX01");
    apply_vector ( 24'b111000111001000010000000,17'b0X1010100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101000010000011  110110100X0XXXX00");
    apply_vector ( 24'b010000110101000010000011,17'b110110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101000010000000  0X1110100X0XXXX00");
    apply_vector ( 24'b111000111101000010000000,17'b0X1110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011000010000000  100001100X0XXXX00");
    apply_vector ( 24'b001000110011000010000000,17'b100001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011000010000001  0X1001100X0XXXX00");
    apply_vector ( 24'b111000111011000010000001,17'b0X1001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111000010000001  110101100X0XXXX00");
    apply_vector ( 24'b010000110111000010000001,17'b110101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111000010000000  0X1101100X0XXXX00");
    apply_vector ( 24'b111000111111000010000000,17'b0X1101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000000010000001  101011000X0XXXX00");
    apply_vector ( 24'b001010110000000010000001,17'b101011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000000010000000  0X0111000X1010011");
    apply_vector ( 24'b111010111000000010000000,17'b0X0111000X1010011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100000010000010  111111000X0010010");
    apply_vector ( 24'b010010110100000010000010,17'b111111000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100000010000001  0X0000100X0010010");
    apply_vector ( 24'b111010111100000010000001,17'b0X0000100X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010000010000000  101000100X0010010");
    apply_vector ( 24'b001010110010000010000000,17'b101000100X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010000010000001  0X0100100X0010010");
    apply_vector ( 24'b111010111010000010000001,17'b0X0100100X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110000010000001  111100100X0010010");
    apply_vector ( 24'b010010110110000010000001,17'b111100100X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110000010000000  0X0010100X0010010");
    apply_vector ( 24'b111010111110000010000000,17'b0X0010100X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001000010000001  101010100X0010010");
    apply_vector ( 24'b001010110001000010000001,17'b101010100X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001000010000000  0X0110100X1110011");
    apply_vector ( 24'b111010111001000010000000,17'b0X0110100X1110011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101000010000011  111110100X0110010");
    apply_vector ( 24'b010010110101000010000011,17'b111110100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101000010000001  0X0001100X0110010");
    apply_vector ( 24'b111010111101000010000001,17'b0X0001100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011000010000000  101001100X0110010");
    apply_vector ( 24'b001010110011000010000000,17'b101001100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011000010000001  0X0101100X0110010");
    apply_vector ( 24'b111010111011000010000001,17'b0X0101100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111000010000001  111101100X0110010");
    apply_vector ( 24'b010010110111000010000001,17'b111101100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111000010000000  0X0011100X0110010");
    apply_vector ( 24'b111010111111000010000000,17'b0X0011100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000000010000001  100111000X0110010");
    apply_vector ( 24'b001001110000000010000001,17'b100111000X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000000010000000  0X1111000X1XXXX01");
    apply_vector ( 24'b111001111000000010000000,17'b0X1111000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100000010000010  110000100X0XXXX00");
    apply_vector ( 24'b010001110100000010000010,17'b110000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100000010000000  0X1000100X0XXXX00");
    apply_vector ( 24'b111001111100000010000000,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010000010000001  100100100X0XXXX00");
    apply_vector ( 24'b001001110010000010000001,17'b100100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010000010000001  0X1100100X0XXXX00");
    apply_vector ( 24'b111001111010000010000001,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110000010000001  110010100X0XXXX00");
    apply_vector ( 24'b010001110110000010000001,17'b110010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110000010000000  0X1010100X0XXXX00");
    apply_vector ( 24'b111001111110000010000000,17'b0X1010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001000010000001  100110100X0XXXX00");
    apply_vector ( 24'b001001110001000010000001,17'b100110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001000010000000  0X1110100X1110011");
    apply_vector ( 24'b111001111001000010000000,17'b0X1110100X1110011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101000010000011  110001100X0110010");
    apply_vector ( 24'b010001110101000010000011,17'b110001100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101000010000000  0X1001100X0110010");
    apply_vector ( 24'b111001111101000010000000,17'b0X1001100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011000010000001  100101100X0110010");
    apply_vector ( 24'b001001110011000010000001,17'b100101100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011000010000001  0X1101100X0110010");
    apply_vector ( 24'b111001111011000010000001,17'b0X1101100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111000010000001  110011100X0110010");
    apply_vector ( 24'b010001110111000010000001,17'b110011100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111000010000000  0X1011100X0110010");
    apply_vector ( 24'b111001111111000010000000,17'b0X1011100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000000010000001  101111000X0110010");
    apply_vector ( 24'b001011110000000010000001,17'b101111000X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000000010000000  0X0000100X1XXXX01");
    apply_vector ( 24'b111011111000000010000000,17'b0X0000100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100000010000010  111000100X0XXXX00");
    apply_vector ( 24'b010011110100000010000010,17'b111000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100000010000001  0X0100100X0XXXX00");
    apply_vector ( 24'b111011111100000010000001,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010000010000001  101100100X0XXXX00");
    apply_vector ( 24'b001011110010000010000001,17'b101100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010000010000001  0X0010100X0XXXX00");
    apply_vector ( 24'b111011111010000010000001,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110000010000001  111010100X0XXXX00");
    apply_vector ( 24'b010011110110000010000001,17'b111010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110000010000000  0X0110100X0XXXX00");
    apply_vector ( 24'b111011111110000010000000,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001000010000001  101110100X0XXXX00");
    apply_vector ( 24'b001011110001000010000001,17'b101110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001000010000000  0X0001100X1110010");
    apply_vector ( 24'b111011111001000010000000,17'b0X0001100X1110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101000010000011  111001100X0110010");
    apply_vector ( 24'b010011110101000010000011,17'b111001100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101000010000001  0X0101100X0110010");
    apply_vector ( 24'b111011111101000010000001,17'b0X0101100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011000010000001  101101100X0110010");
    apply_vector ( 24'b001011110011000010000001,17'b101101100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011000010000001  0X0011100X0110010");
    apply_vector ( 24'b111011111011000010000001,17'b0X0011100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111000010000001  111011100X0110010");
    apply_vector ( 24'b010011110111000010000001,17'b111011100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111000010000000  0X0111100X0110010");
    apply_vector ( 24'b111011111111000010000000,17'b0X0111100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000000010000001  101000000X0110010");
    apply_vector ( 24'b001100000000000010000001,17'b101000000X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000000010000000  0X0100000X1110011");
    apply_vector ( 24'b111100001000000010000000,17'b0X0100000X1110011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100000010000010  111100000X0110010");
    apply_vector ( 24'b010100000100000010000010,17'b111100000X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100000010000000  0X0010000X0110010");
    apply_vector ( 24'b111100001100000010000000,17'b0X0010000X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010000010000000  101010000X0110010");
    apply_vector ( 24'b001100000010000010000000,17'b101010000X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010000010000000  0X0110000X0110010");
    apply_vector ( 24'b111100001010000010000000,17'b0X0110000X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110000010000000  111110000X0110010");
    apply_vector ( 24'b010100000110000010000000,17'b111110000X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110000010000001  0X0001000X0110010");
    apply_vector ( 24'b111100001110000010000001,17'b0X0001000X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001000010000001  101001000X0110010");
    apply_vector ( 24'b001100000001000010000001,17'b101001000X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001000010000000  0X0101000X1001011");
    apply_vector ( 24'b111100001001000010000000,17'b0X0101000X1001011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101000010000011  111101000X0001010");
    apply_vector ( 24'b010100000101000010000011,17'b111101000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101000010000000  0X0011000X0001010");
    apply_vector ( 24'b111100001101000010000000,17'b0X0011000X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011000010000000  101011000X0001010");
    apply_vector ( 24'b001100000011000010000000,17'b101011000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011000010000000  0X0111000X0001010");
    apply_vector ( 24'b111100001011000010000000,17'b0X0111000X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111000010000000  111111000X0001010");
    apply_vector ( 24'b010100000111000010000000,17'b111111000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111000010000001  0X0000100X0001010");
    apply_vector ( 24'b111100001111000010000001,17'b0X0000100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000000010000001  100100000X0001010");
    apply_vector ( 24'b001110000000000010000001,17'b100100000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000000010000000  0X1100000X1XXXX01");
    apply_vector ( 24'b111110001000000010000000,17'b0X1100000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100000010000010  110010000X0XXXX00");
    apply_vector ( 24'b010110000100000010000010,17'b110010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100000010000001  0X1010000X0XXXX00");
    apply_vector ( 24'b111110001100000010000001,17'b0X1010000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010000010000000  100110000X0XXXX00");
    apply_vector ( 24'b001110000010000010000000,17'b100110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010000010000000  0X1110000X0XXXX00");
    apply_vector ( 24'b111110001010000010000000,17'b0X1110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110000010000000  110001000X0XXXX00");
    apply_vector ( 24'b010110000110000010000000,17'b110001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110000010000001  0X1001000X0XXXX00");
    apply_vector ( 24'b111110001110000010000001,17'b0X1001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001000010000001  100101000X0XXXX00");
    apply_vector ( 24'b001110000001000010000001,17'b100101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001000010000000  0X1101000X1XXXX01");
    apply_vector ( 24'b111110001001000010000000,17'b0X1101000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101000010000011  110011000X0XXXX00");
    apply_vector ( 24'b010110000101000010000011,17'b110011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101000010000001  0X1011000X0XXXX00");
    apply_vector ( 24'b111110001101000010000001,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011000010000000  100111000X0XXXX00");
    apply_vector ( 24'b001110000011000010000000,17'b100111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111110001011000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111000010000000  110000100X0XXXX00");
    apply_vector ( 24'b010110000111000010000000,17'b110000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111000010000001  0X1000100X0XXXX00");
    apply_vector ( 24'b111110001111000010000001,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000000010000001  101100000X0XXXX00");
    apply_vector ( 24'b001101000000000010000001,17'b101100000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101001000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000000010000000  0X0010000X1101011");
    apply_vector ( 24'b111101001000000010000000,17'b0X0010000X1101011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100000010000010  111010000X0101010");
    apply_vector ( 24'b010101000100000010000010,17'b111010000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100000010000000  0X0110000X0101010");
    apply_vector ( 24'b111101001100000010000000,17'b0X0110000X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010000010000001  101110000X0101010");
    apply_vector ( 24'b001101000010000010000001,17'b101110000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010000010000000  0X0001000X0101010");
    apply_vector ( 24'b111101001010000010000000,17'b0X0001000X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110000010000000  111001000X0101010");
    apply_vector ( 24'b010101000110000010000000,17'b111001000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110000010000001  0X0101000X0101010");
    apply_vector ( 24'b111101001110000010000001,17'b0X0101000X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001000010000001  101101000X0101010");
    apply_vector ( 24'b001101000001000010000001,17'b101101000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001000010000000  0X0011000X1001010");
    apply_vector ( 24'b111101001001000010000000,17'b0X0011000X1001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101000010000011  111011000X0001010");
    apply_vector ( 24'b010101000101000010000011,17'b111011000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101000010000000  0X0111000X0001010");
    apply_vector ( 24'b111101001101000010000000,17'b0X0111000X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011000010000001  101111000X0001010");
    apply_vector ( 24'b001101000011000010000001,17'b101111000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011000010000000  0X0000100X0001010");
    apply_vector ( 24'b111101001011000010000000,17'b0X0000100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111000010000000  111000100X0001010");
    apply_vector ( 24'b010101000111000010000000,17'b111000100X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111000010000001  0X0100100X0001010");
    apply_vector ( 24'b111101001111000010000001,17'b0X0100100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000000010000001  100010000X0001010");
    apply_vector ( 24'b001111000000000010000001,17'b100010000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000000010000000  0X1010000X1001011");
    apply_vector ( 24'b111111001000000010000000,17'b0X1010000X1001011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100000010000010  110110000X0001010");
    apply_vector ( 24'b010111000100000010000010,17'b110110000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100000010000001  0X1110000X0001010");
    apply_vector ( 24'b111111001100000010000001,17'b0X1110000X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010000010000001  100001000X0001010");
    apply_vector ( 24'b001111000010000010000001,17'b100001000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010000010000000  0X1001000X0001010");
    apply_vector ( 24'b111111001010000010000000,17'b0X1001000X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110000010000000  110101000X0001010");
    apply_vector ( 24'b010111000110000010000000,17'b110101000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110000010000001  0X1101000X0001010");
    apply_vector ( 24'b111111001110000010000001,17'b0X1101000X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001000010000001  100011000X0001010");
    apply_vector ( 24'b001111000001000010000001,17'b100011000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001000010000000  0X1011000X1001011");
    apply_vector ( 24'b111111001001000010000000,17'b0X1011000X1001011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101000010000011  110111000X0001010");
    apply_vector ( 24'b010111000101000010000011,17'b110111000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101000010000001  0X1111000X0001010");
    apply_vector ( 24'b111111001101000010000001,17'b0X1111000X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011000010000001  100000100X0001010");
    apply_vector ( 24'b001111000011000010000001,17'b100000100X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011000010000000  0X1000100X0001010");
    apply_vector ( 24'b111111001011000010000000,17'b0X1000100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111000010000000  110100100X0001010");
    apply_vector ( 24'b010111000111000010000000,17'b110100100X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111000010000001  0X1100100X0001010");
    apply_vector ( 24'b111111001111000010000001,17'b0X1100100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000000010000001  101010000X0001010");
    apply_vector ( 24'b001100100000000010000001,17'b101010000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000000010000000  0X0110000X1XXXX01");
    apply_vector ( 24'b111100101000000010000000,17'b0X0110000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100000010000010  111110000X0XXXX00");
    apply_vector ( 24'b010100100100000010000010,17'b111110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100000010000000  0X0001000X0XXXX00");
    apply_vector ( 24'b111100101100000010000000,17'b0X0001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010000010000000  101001000X0XXXX00");
    apply_vector ( 24'b001100100010000010000000,17'b101001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010000010000001  0X0101000X0XXXX00");
    apply_vector ( 24'b111100101010000010000001,17'b0X0101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110000010000000  111101000X0XXXX00");
    apply_vector ( 24'b010100100110000010000000,17'b111101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110000010000001  0X0011000X0XXXX00");
    apply_vector ( 24'b111100101110000010000001,17'b0X0011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001000010000001  101011000X0XXXX00");
    apply_vector ( 24'b001100100001000010000001,17'b101011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001000010000000  0X0111000X1XXXX01");
    apply_vector ( 24'b111100101001000010000000,17'b0X0111000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101000010000011  111111000X0XXXX00");
    apply_vector ( 24'b010100100101000010000011,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101000010000000  0X0000100X0XXXX00");
    apply_vector ( 24'b111100101101000010000000,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011000010000000  101000100X0XXXX00");
    apply_vector ( 24'b001100100011000010000000,17'b101000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011000010000001  0X0100100X0XXXX00");
    apply_vector ( 24'b111100101011000010000001,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111000010000000  111100100X0XXXX00");
    apply_vector ( 24'b010100100111000010000000,17'b111100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111000010000001  0X0010100X0XXXX00");
    apply_vector ( 24'b111100101111000010000001,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000000010000001  100110000X0XXXX00");
    apply_vector ( 24'b001110100000000010000001,17'b100110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110101000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000000010000000  0X1110000X1010011");
    apply_vector ( 24'b111110101000000010000000,17'b0X1110000X1010011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100000010000010  110001000X0010010");
    apply_vector ( 24'b010110100100000010000010,17'b110001000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100000010000001  0X1001000X0010010");
    apply_vector ( 24'b111110101100000010000001,17'b0X1001000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010000010000000  100101000X0010010");
    apply_vector ( 24'b001110100010000010000000,17'b100101000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010000010000001  0X1101000X0010010");
    apply_vector ( 24'b111110101010000010000001,17'b0X1101000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110000010000000  110011000X0010010");
    apply_vector ( 24'b010110100110000010000000,17'b110011000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110000010000001  0X1011000X0010010");
    apply_vector ( 24'b111110101110000010000001,17'b0X1011000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001000010000001  100111000X0010010");
    apply_vector ( 24'b001110100001000010000001,17'b100111000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001000010000000  0X1111000X1111111");
    apply_vector ( 24'b111110101001000010000000,17'b0X1111000X1111111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101000010000011  110000100X0111110");
    apply_vector ( 24'b010110100101000010000011,17'b110000100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101000010000001  0X1000100X0111110");
    apply_vector ( 24'b111110101101000010000001,17'b0X1000100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011000010000000  100100100X0111110");
    apply_vector ( 24'b001110100011000010000000,17'b100100100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011000010000001  0X1100100X0111110");
    apply_vector ( 24'b111110101011000010000001,17'b0X1100100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111000010000000  110010100X0111110");
    apply_vector ( 24'b010110100111000010000000,17'b110010100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111000010000001  0X1010100X0111110");
    apply_vector ( 24'b111110101111000010000001,17'b0X1010100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000000010000001  101110000X0111110");
    apply_vector ( 24'b001101100000000010000001,17'b101110000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000000010000000  0X0001000X1XXXX01");
    apply_vector ( 24'b111101101000000010000000,17'b0X0001000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100000010000010  111001000X0XXXX00");
    apply_vector ( 24'b010101100100000010000010,17'b111001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100000010000000  0X0101000X0XXXX00");
    apply_vector ( 24'b111101101100000010000000,17'b0X0101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010000010000001  101101000X0XXXX00");
    apply_vector ( 24'b001101100010000010000001,17'b101101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010000010000001  0X0011000X0XXXX00");
    apply_vector ( 24'b111101101010000010000001,17'b0X0011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110000010000000  111011000X0XXXX00");
    apply_vector ( 24'b010101100110000010000000,17'b111011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110000010000001  0X0111000X0XXXX00");
    apply_vector ( 24'b111101101110000010000001,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001000010000001  101111000X0XXXX00");
    apply_vector ( 24'b001101100001000010000001,17'b101111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001000010000000  0X0000100X1001011");
    apply_vector ( 24'b111101101001000010000000,17'b0X0000100X1001011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101000010000011  111000100X0001010");
    apply_vector ( 24'b010101100101000010000011,17'b111000100X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101000010000000  0X0100100X0001010");
    apply_vector ( 24'b111101101101000010000000,17'b0X0100100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011000010000001  101100100X0001010");
    apply_vector ( 24'b001101100011000010000001,17'b101100100X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011000010000001  0X0010100X0001010");
    apply_vector ( 24'b111101101011000010000001,17'b0X0010100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111000010000000  111010100X0001010");
    apply_vector ( 24'b010101100111000010000000,17'b111010100X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111000010000001  0X0110100X0001010");
    apply_vector ( 24'b111101101111000010000001,17'b0X0110100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000000010000001  100001000X0001010");
    apply_vector ( 24'b001111100000000010000001,17'b100001000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000000010000000  0X1001000X1XXXX01");
    apply_vector ( 24'b111111101000000010000000,17'b0X1001000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100000010000010  110101000X0XXXX00");
    apply_vector ( 24'b010111100100000010000010,17'b110101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100000010000001  0X1101000X0XXXX00");
    apply_vector ( 24'b111111101100000010000001,17'b0X1101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010000010000001  100011000X0XXXX00");
    apply_vector ( 24'b001111100010000010000001,17'b100011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010000010000001  0X1011000X0XXXX00");
    apply_vector ( 24'b111111101010000010000001,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110000010000000  110111000X0XXXX00");
    apply_vector ( 24'b010111100110000010000000,17'b110111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110000010000001  0X1111000X0XXXX00");
    apply_vector ( 24'b111111101110000010000001,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001000010000001  100000100X0XXXX00");
    apply_vector ( 24'b001111100001000010000001,17'b100000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001000010000000  0X1000100X1XXXX01");
    apply_vector ( 24'b111111101001000010000000,17'b0X1000100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101000010000011  110100100X0XXXX00");
    apply_vector ( 24'b010111100101000010000011,17'b110100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101000010000001  0X1100100X0XXXX00");
    apply_vector ( 24'b111111101101000010000001,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011000010000001  100010100X0XXXX00");
    apply_vector ( 24'b001111100011000010000001,17'b100010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011000010000001  0X1010100X0XXXX00");
    apply_vector ( 24'b111111101011000010000001,17'b0X1010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111000010000000  110110100X0XXXX00");
    apply_vector ( 24'b010111100111000010000000,17'b110110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111000010000001  0X1110100X0XXXX00");
    apply_vector ( 24'b111111101111000010000001,17'b0X1110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000000010000001  101001000X0XXXX00");
    apply_vector ( 24'b001100010000000010000001,17'b101001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000000010000000  0X0101000X1111011");
    apply_vector ( 24'b111100011000000010000000,17'b0X0101000X1111011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100000010000010  111101000X0111010");
    apply_vector ( 24'b010100010100000010000010,17'b111101000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100000010000000  0X0011000X0111010");
    apply_vector ( 24'b111100011100000010000000,17'b0X0011000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010000010000000  101011000X0111010");
    apply_vector ( 24'b001100010010000010000000,17'b101011000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010000010000000  0X0111000X0111010");
    apply_vector ( 24'b111100011010000010000000,17'b0X0111000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110000010000001  111111000X0111010");
    apply_vector ( 24'b010100010110000010000001,17'b111111000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110000010000001  0X0000100X0111010");
    apply_vector ( 24'b111100011110000010000001,17'b0X0000100X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001000010000001  101000100X0111010");
    apply_vector ( 24'b001100010001000010000001,17'b101000100X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001000010000000  0X0100100X1XXXX01");
    apply_vector ( 24'b111100011001000010000000,17'b0X0100100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101000010000011  111100100X0XXXX00");
    apply_vector ( 24'b010100010101000010000011,17'b111100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101000010000000  0X0010100X0XXXX00");
    apply_vector ( 24'b111100011101000010000000,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011000010000000  101010100X0XXXX00");
    apply_vector ( 24'b001100010011000010000000,17'b101010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011000010000000  0X0110100X0XXXX00");
    apply_vector ( 24'b111100011011000010000000,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111000010000001  111110100X0XXXX00");
    apply_vector ( 24'b010100010111000010000001,17'b111110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111000010000001  0X0001100X0XXXX00");
    apply_vector ( 24'b111100011111000010000001,17'b0X0001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000000010000001  100101000X0XXXX00");
    apply_vector ( 24'b001110010000000010000001,17'b100101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000000010000000  0X1101000X1101011");
    apply_vector ( 24'b111110011000000010000000,17'b0X1101000X1101011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100000010000010  110011000X0101010");
    apply_vector ( 24'b010110010100000010000010,17'b110011000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100000010000001  0X1011000X0101010");
    apply_vector ( 24'b111110011100000010000001,17'b0X1011000X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010000010000000  100111000X0101010");
    apply_vector ( 24'b001110010010000010000000,17'b100111000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010000010000000  0X1111000X0101010");
    apply_vector ( 24'b111110011010000010000000,17'b0X1111000X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110000010000001  110000100X0101010");
    apply_vector ( 24'b010110010110000010000001,17'b110000100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110000010000001  0X1000100X0101010");
    apply_vector ( 24'b111110011110000010000001,17'b0X1000100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001000010000001  100100100X0101010");
    apply_vector ( 24'b001110010001000010000001,17'b100100100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001000010000000  0X1100100X1101011");
    apply_vector ( 24'b111110011001000010000000,17'b0X1100100X1101011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101000010000011  110010100X0101010");
    apply_vector ( 24'b010110010101000010000011,17'b110010100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101000010000001  0X1010100X0101010");
    apply_vector ( 24'b111110011101000010000001,17'b0X1010100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011000010000000  100110100X0101010");
    apply_vector ( 24'b001110010011000010000000,17'b100110100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011000010000000  0X1110100X0101010");
    apply_vector ( 24'b111110011011000010000000,17'b0X1110100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111000010000001  110001100X0101010");
    apply_vector ( 24'b010110010111000010000001,17'b110001100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111000010000001  0X1001100X0101010");
    apply_vector ( 24'b111110011111000010000001,17'b0X1001100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000000010000001  101101000X0101010");
    apply_vector ( 24'b001101010000000010000001,17'b101101000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000000010000000  0X0011000X1101010");
    apply_vector ( 24'b111101011000000010000000,17'b0X0011000X1101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100000010000010  111011000X0101010");
    apply_vector ( 24'b010101010100000010000010,17'b111011000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100000010000000  0X0111000X0101010");
    apply_vector ( 24'b111101011100000010000000,17'b0X0111000X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010000010000001  101111000X0101010");
    apply_vector ( 24'b001101010010000010000001,17'b101111000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010000010000000  0X0000100X0101010");
    apply_vector ( 24'b111101011010000010000000,17'b0X0000100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110000010000001  111000100X0101010");
    apply_vector ( 24'b010101010110000010000001,17'b111000100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110000010000001  0X0100100X0101010");
    apply_vector ( 24'b111101011110000010000001,17'b0X0100100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001000010000001  101100100X0101010");
    apply_vector ( 24'b001101010001000010000001,17'b101100100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001000010000000  0X0010100X1001011");
    apply_vector ( 24'b111101011001000010000000,17'b0X0010100X1001011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101000010000011  111010100X0001010");
    apply_vector ( 24'b010101010101000010000011,17'b111010100X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101000010000000  0X0110100X0001010");
    apply_vector ( 24'b111101011101000010000000,17'b0X0110100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011000010000001  101110100X0001010");
    apply_vector ( 24'b001101010011000010000001,17'b101110100X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011000010000000  0X0001100X0001010");
    apply_vector ( 24'b111101011011000010000000,17'b0X0001100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111000010000001  111001100X0001010");
    apply_vector ( 24'b010101010111000010000001,17'b111001100X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111000010000001  0X0101100X0001010");
    apply_vector ( 24'b111101011111000010000001,17'b0X0101100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000000010000001  100011000X0001010");
    apply_vector ( 24'b001111010000000010000001,17'b100011000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000000010000000  0X1011000X1XXXX01");
    apply_vector ( 24'b111111011000000010000000,17'b0X1011000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100000010000010  110111000X0XXXX00");
    apply_vector ( 24'b010111010100000010000010,17'b110111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100000010000001  0X1111000X0XXXX00");
    apply_vector ( 24'b111111011100000010000001,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010000010000001  100000100X0XXXX00");
    apply_vector ( 24'b001111010010000010000001,17'b100000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010000010000000  0X1000100X0XXXX00");
    apply_vector ( 24'b111111011010000010000000,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110000010000001  110100100X0XXXX00");
    apply_vector ( 24'b010111010110000010000001,17'b110100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110000010000001  0X1100100X0XXXX00");
    apply_vector ( 24'b111111011110000010000001,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001000010000001  100010100X0XXXX00");
    apply_vector ( 24'b001111010001000010000001,17'b100010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111011001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001000010000000  0X1010100X1XXXX01");
    apply_vector ( 24'b111111011001000010000000,17'b0X1010100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101000010000011  110110100X0XXXX00");
    apply_vector ( 24'b010111010101000010000011,17'b110110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101000010000001  0X1110100X0XXXX00");
    apply_vector ( 24'b111111011101000010000001,17'b0X1110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011000010000001  100001100X0XXXX00");
    apply_vector ( 24'b001111010011000010000001,17'b100001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011000010000000  0X1001100X0XXXX00");
    apply_vector ( 24'b111111011011000010000000,17'b0X1001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111000010000001  110101100X0XXXX00");
    apply_vector ( 24'b010111010111000010000001,17'b110101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111000010000001  0X1101100X0XXXX00");
    apply_vector ( 24'b111111011111000010000001,17'b0X1101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000000010000001  101011000X0XXXX00");
    apply_vector ( 24'b001100110000000010000001,17'b101011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000000010000000  0X0111000X1101011");
    apply_vector ( 24'b111100111000000010000000,17'b0X0111000X1101011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100000010000010  111111000X0101010");
    apply_vector ( 24'b010100110100000010000010,17'b111111000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100000010000000  0X0000100X0101010");
    apply_vector ( 24'b111100111100000010000000,17'b0X0000100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010000010000000  101000100X0101010");
    apply_vector ( 24'b001100110010000010000000,17'b101000100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010000010000001  0X0100100X0101010");
    apply_vector ( 24'b111100111010000010000001,17'b0X0100100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110000010000001  111100100X0101010");
    apply_vector ( 24'b010100110110000010000001,17'b111100100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110000010000001  0X0010100X0101010");
    apply_vector ( 24'b111100111110000010000001,17'b0X0010100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001000010000001  101010100X0101010");
    apply_vector ( 24'b001100110001000010000001,17'b101010100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001000010000000  0X0110100X1011011");
    apply_vector ( 24'b111100111001000010000000,17'b0X0110100X1011011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101000010000011  111110100X0011010");
    apply_vector ( 24'b010100110101000010000011,17'b111110100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101000010000000  0X0001100X0011010");
    apply_vector ( 24'b111100111101000010000000,17'b0X0001100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011000010000000  101001100X0011010");
    apply_vector ( 24'b001100110011000010000000,17'b101001100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011000010000001  0X0101100X0011010");
    apply_vector ( 24'b111100111011000010000001,17'b0X0101100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111000010000001  111101100X0011010");
    apply_vector ( 24'b010100110111000010000001,17'b111101100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111000010000001  0X0011100X0011010");
    apply_vector ( 24'b111100111111000010000001,17'b0X0011100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000000010000001  100111000X0011010");
    apply_vector ( 24'b001110110000000010000001,17'b100111000X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000000010000000  0X1111000X1XXXX01");
    apply_vector ( 24'b111110111000000010000000,17'b0X1111000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100000010000010  110000100X0XXXX00");
    apply_vector ( 24'b010110110100000010000010,17'b110000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100000010000001  0X1000100X0XXXX00");
    apply_vector ( 24'b111110111100000010000001,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010000010000000  100100100X0XXXX00");
    apply_vector ( 24'b001110110010000010000000,17'b100100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010000010000001  0X1100100X0XXXX00");
    apply_vector ( 24'b111110111010000010000001,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110000010000001  110010100X0XXXX00");
    apply_vector ( 24'b010110110110000010000001,17'b110010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110000010000001  0X1010100X0XXXX00");
    apply_vector ( 24'b111110111110000010000001,17'b0X1010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001000010000001  100110100X0XXXX00");
    apply_vector ( 24'b001110110001000010000001,17'b100110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001000010000000  0X1110100X1XXXX01");
    apply_vector ( 24'b111110111001000010000000,17'b0X1110100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101000010000011  110001100X0XXXX00");
    apply_vector ( 24'b010110110101000010000011,17'b110001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101000010000001  0X1001100X0XXXX00");
    apply_vector ( 24'b111110111101000010000001,17'b0X1001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011000010000000  100101100X0XXXX00");
    apply_vector ( 24'b001110110011000010000000,17'b100101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011000010000001  0X1101100X0XXXX00");
    apply_vector ( 24'b111110111011000010000001,17'b0X1101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111000010000001  110011100X0XXXX00");
    apply_vector ( 24'b010110110111000010000001,17'b110011100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111000010000001  0X1011100X0XXXX00");
    apply_vector ( 24'b111110111111000010000001,17'b0X1011100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000000010000001  101111000X0XXXX00");
    apply_vector ( 24'b001101110000000010000001,17'b101111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000000010000000  0X0000100X1101011");
    apply_vector ( 24'b111101111000000010000000,17'b0X0000100X1101011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100000010000010  111000100X0101010");
    apply_vector ( 24'b010101110100000010000010,17'b111000100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100000010000000  0X0100100X0101010");
    apply_vector ( 24'b111101111100000010000000,17'b0X0100100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010000010000001  101100100X0101010");
    apply_vector ( 24'b001101110010000010000001,17'b101100100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010000010000001  0X0010100X0101010");
    apply_vector ( 24'b111101111010000010000001,17'b0X0010100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110000010000001  111010100X0101010");
    apply_vector ( 24'b010101110110000010000001,17'b111010100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110000010000001  0X0110100X0101010");
    apply_vector ( 24'b111101111110000010000001,17'b0X0110100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001000010000001  101110100X0101010");
    apply_vector ( 24'b001101110001000010000001,17'b101110100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001000010000000  0X0001100X1XXXX01");
    apply_vector ( 24'b111101111001000010000000,17'b0X0001100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101000010000011  111001100X0XXXX00");
    apply_vector ( 24'b010101110101000010000011,17'b111001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101000010000000  0X0101100X0XXXX00");
    apply_vector ( 24'b111101111101000010000000,17'b0X0101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011000010000001  101101100X0XXXX00");
    apply_vector ( 24'b001101110011000010000001,17'b101101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011000010000001  0X0011100X0XXXX00");
    apply_vector ( 24'b111101111011000010000001,17'b0X0011100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111000010000001  111011100X0XXXX00");
    apply_vector ( 24'b010101110111000010000001,17'b111011100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111000010000001  0X0111100X0XXXX00");
    apply_vector ( 24'b111101111111000010000001,17'b0X0111100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000000010000001  100000100X0XXXX00");
    apply_vector ( 24'b001111110000000010000001,17'b100000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111111000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000000010000000  0X1000100X1011111");
    apply_vector ( 24'b111111111000000010000000,17'b0X1000100X1011111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100000010000010  110100100X0011110");
    apply_vector ( 24'b010111110100000010000010,17'b110100100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100000010000001  0X1100100X0011110");
    apply_vector ( 24'b111111111100000010000001,17'b0X1100100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010000010000001  100010100X0011110");
    apply_vector ( 24'b001111110010000010000001,17'b100010100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010000010000001  0X1010100X0011110");
    apply_vector ( 24'b111111111010000010000001,17'b0X1010100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110000010000001  110110100X0011110");
    apply_vector ( 24'b010111110110000010000001,17'b110110100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110000010000001  0X1110100X0011110");
    apply_vector ( 24'b111111111110000010000001,17'b0X1110100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001000010000001  100001100X0011110");
    apply_vector ( 24'b001111110001000010000001,17'b100001100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001000010000000  0X1001100X1110011");
    apply_vector ( 24'b111111111001000010000000,17'b0X1001100X1110011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101000010000011  110101100X0110010");
    apply_vector ( 24'b010111110101000010000011,17'b110101100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101000010000001  0X1101100X0110010");
    apply_vector ( 24'b111111111101000010000001,17'b0X1101100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011000010000001  100011100X0110010");
    apply_vector ( 24'b001111110011000010000001,17'b100011100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011000010000001  0X1011100X0110010");
    apply_vector ( 24'b111111111011000010000001,17'b0X1011100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111000010000001  110111100X0110010");
    apply_vector ( 24'b010111110111000010000001,17'b110111100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111000010000001  0X1111100X0110010");
    apply_vector ( 24'b111111111111000010000001,17'b0X1111100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000000010000001  100000000X0110010");
    apply_vector ( 24'b001000000000000010000001,17'b100000000X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000001000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000000010000000  0X1000000X1XXXX01");
    apply_vector ( 24'b111000001000000010000000,17'b0X1000000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100000010000010  110100000X0XXXX00");
    apply_vector ( 24'b010000000100000010000010,17'b110100000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100000010000000  0X1100000X0XXXX00");
    apply_vector ( 24'b111000001100000010000000,17'b0X1100000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010000010000000  100010000X0XXXX00");
    apply_vector ( 24'b001000000010000010000000,17'b100010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010000010000000  0X1010000X0XXXX00");
    apply_vector ( 24'b111000001010000010000000,17'b0X1010000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110000010000000  110110000X0XXXX00");
    apply_vector ( 24'b010000000110000010000000,17'b110110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110000010000000  0X1110000X0XXXX00");
    apply_vector ( 24'b111000001110000010000000,17'b0X1110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001000010000000  100001000X0XXXX00");
    apply_vector ( 24'b001000000001000010000000,17'b100001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001000010000001  0X1001000X1XXXX01");
    apply_vector ( 24'b111000001001000010000001,17'b0X1001000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101000010000011  110101000X0XXXX00");
    apply_vector ( 24'b010000000101000010000011,17'b110101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101000010000000  0X1101000X0XXXX00");
    apply_vector ( 24'b111000001101000010000000,17'b0X1101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011000010000000  100011000X0XXXX00");
    apply_vector ( 24'b001000000011000010000000,17'b100011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011000010000000  0X1011000X0XXXX00");
    apply_vector ( 24'b111000001011000010000000,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111000010000000  110111000X0XXXX00");
    apply_vector ( 24'b010000000111000010000000,17'b110111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111000001111000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010000000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000000010000000  101000000X0XXXX00");
    apply_vector ( 24'b001010000000000010000000,17'b101000000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000000010000001  0X0100000X1001111");
    apply_vector ( 24'b111010001000000010000001,17'b0X0100000X1001111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100000010000010  111100000X0001110");
    apply_vector ( 24'b010010000100000010000010,17'b111100000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100000010000001  0X0010000X0001110");
    apply_vector ( 24'b111010001100000010000001,17'b0X0010000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010000010000000  101010000X0001110");
    apply_vector ( 24'b001010000010000010000000,17'b101010000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010000010000000  0X0110000X0001110");
    apply_vector ( 24'b111010001010000010000000,17'b0X0110000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110000010000000  111110000X0001110");
    apply_vector ( 24'b010010000110000010000000,17'b111110000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110000010000000  0X0001000X0001110");
    apply_vector ( 24'b111010001110000010000000,17'b0X0001000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001000010000000  101001000X0001110");
    apply_vector ( 24'b001010000001000010000000,17'b101001000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001000010000001  0X0101000X1100011");
    apply_vector ( 24'b111010001001000010000001,17'b0X0101000X1100011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101000010000011  111101000X0100010");
    apply_vector ( 24'b010010000101000010000011,17'b111101000X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101000010000001  0X0011000X0100010");
    apply_vector ( 24'b111010001101000010000001,17'b0X0011000X0100010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011000010000000  101011000X0100010");
    apply_vector ( 24'b001010000011000010000000,17'b101011000X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011000010000000  0X0111000X0100010");
    apply_vector ( 24'b111010001011000010000000,17'b0X0111000X0100010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111000010000000  111111000X0100010");
    apply_vector ( 24'b010010000111000010000000,17'b111111000X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111000010000000  0X0000100X0100010");
    apply_vector ( 24'b111010001111000010000000,17'b0X0000100X0100010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001000000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000000010000000  100100000X0100010");
    apply_vector ( 24'b001001000000000010000000,17'b100100000X0100010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000000010000001  0X1100000X1XXXX01");
    apply_vector ( 24'b111001001000000010000001,17'b0X1100000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100000010000010  110010000X0XXXX00");
    apply_vector ( 24'b010001000100000010000010,17'b110010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100000010000000  0X1010000X0XXXX00");
    apply_vector ( 24'b111001001100000010000000,17'b0X1010000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010000010000001  100110000X0XXXX00");
    apply_vector ( 24'b001001000010000010000001,17'b100110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010000010000000  0X1110000X0XXXX00");
    apply_vector ( 24'b111001001010000010000000,17'b0X1110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110000010000000  110001000X0XXXX00");
    apply_vector ( 24'b010001000110000010000000,17'b110001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110000010000000  0X1001000X0XXXX00");
    apply_vector ( 24'b111001001110000010000000,17'b0X1001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001000010000000  100101000X0XXXX00");
    apply_vector ( 24'b001001000001000010000000,17'b100101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001000010000001  0X1101000X1010111");
    apply_vector ( 24'b111001001001000010000001,17'b0X1101000X1010111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101000010000011  110011000X0010110");
    apply_vector ( 24'b010001000101000010000011,17'b110011000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101000010000000  0X1011000X0010110");
    apply_vector ( 24'b111001001101000010000000,17'b0X1011000X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011000010000001  100111000X0010110");
    apply_vector ( 24'b001001000011000010000001,17'b100111000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011000010000000  0X1111000X0010110");
    apply_vector ( 24'b111001001011000010000000,17'b0X1111000X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111000010000000  110000100X0010110");
    apply_vector ( 24'b010001000111000010000000,17'b110000100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001001111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111000010000000  0X1000100X0010110");
    apply_vector ( 24'b111001001111000010000000,17'b0X1000100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011000000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000000010000000  101100000X0010110");
    apply_vector ( 24'b001011000000000010000000,17'b101100000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000000010000001  0X0010000X1XXXX01");
    apply_vector ( 24'b111011001000000010000001,17'b0X0010000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100000010000010  111010000X0XXXX00");
    apply_vector ( 24'b010011000100000010000010,17'b111010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100000010000001  0X0110000X0XXXX00");
    apply_vector ( 24'b111011001100000010000001,17'b0X0110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010000010000001  101110000X0XXXX00");
    apply_vector ( 24'b001011000010000010000001,17'b101110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010000010000000  0X0001000X0XXXX00");
    apply_vector ( 24'b111011001010000010000000,17'b0X0001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110000010000000  111001000X0XXXX00");
    apply_vector ( 24'b010011000110000010000000,17'b111001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110000010000000  0X0101000X0XXXX00");
    apply_vector ( 24'b111011001110000010000000,17'b0X0101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001000010000000  101101000X0XXXX00");
    apply_vector ( 24'b001011000001000010000000,17'b101101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001000010000001  0X0011000X1XXXX01");
    apply_vector ( 24'b111011001001000010000001,17'b0X0011000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101000010000011  111011000X0XXXX00");
    apply_vector ( 24'b010011000101000010000011,17'b111011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101000010000001  0X0111000X0XXXX00");
    apply_vector ( 24'b111011001101000010000001,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011000010000001  101111000X0XXXX00");
    apply_vector ( 24'b001011000011000010000001,17'b101111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011000010000000  0X0000100X0XXXX00");
    apply_vector ( 24'b111011001011000010000000,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111000010000000  111000100X0XXXX00");
    apply_vector ( 24'b010011000111000010000000,17'b111000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111000010000000  0X0100100X0XXXX00");
    apply_vector ( 24'b111011001111000010000000,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000100000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000000010000000  100010000X0XXXX00");
    apply_vector ( 24'b001000100000000010000000,17'b100010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000000010000001  0X1010000X1100111");
    apply_vector ( 24'b111000101000000010000001,17'b0X1010000X1100111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100000010000010  110110000X0100110");
    apply_vector ( 24'b010000100100000010000010,17'b110110000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100000010000000  0X1110000X0100110");
    apply_vector ( 24'b111000101100000010000000,17'b0X1110000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010000010000000  100001000X0100110");
    apply_vector ( 24'b001000100010000010000000,17'b100001000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010000010000001  0X1001000X0100110");
    apply_vector ( 24'b111000101010000010000001,17'b0X1001000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110000010000000  110101000X0100110");
    apply_vector ( 24'b010000100110000010000000,17'b110101000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110000010000000  0X1101000X0100110");
    apply_vector ( 24'b111000101110000010000000,17'b0X1101000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000100001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001000010000000  100011000X0100110");
    apply_vector ( 24'b001000100001000010000000,17'b100011000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001000010000001  0X1011000X1010111");
    apply_vector ( 24'b111000101001000010000001,17'b0X1011000X1010111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101000010000011  110111000X0010110");
    apply_vector ( 24'b010000100101000010000011,17'b110111000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101000010000000  0X1111000X0010110");
    apply_vector ( 24'b111000101101000010000000,17'b0X1111000X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011000010000000  100000100X0010110");
    apply_vector ( 24'b001000100011000010000000,17'b100000100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011000010000001  0X1000100X0010110");
    apply_vector ( 24'b111000101011000010000001,17'b0X1000100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111000010000000  110100100X0010110");
    apply_vector ( 24'b010000100111000010000000,17'b110100100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111000010000000  0X1100100X0010110");
    apply_vector ( 24'b111000101111000010000000,17'b0X1100100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010100000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000000010000000  101010000X0010110");
    apply_vector ( 24'b001010100000000010000000,17'b101010000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000000010000001  0X0110000X1XXXX01");
    apply_vector ( 24'b111010101000000010000001,17'b0X0110000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100000010000010  111110000X0XXXX00");
    apply_vector ( 24'b010010100100000010000010,17'b111110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100000010000001  0X0001000X0XXXX00");
    apply_vector ( 24'b111010101100000010000001,17'b0X0001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010000010000000  101001000X0XXXX00");
    apply_vector ( 24'b001010100010000010000000,17'b101001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010000010000001  0X0101000X0XXXX00");
    apply_vector ( 24'b111010101010000010000001,17'b0X0101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110000010000000  111101000X0XXXX00");
    apply_vector ( 24'b010010100110000010000000,17'b111101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010101110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110000010000000  0X0011000X0XXXX00");
    apply_vector ( 24'b111010101110000010000000,17'b0X0011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010100001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001000010000000  101011000X0XXXX00");
    apply_vector ( 24'b001010100001000010000000,17'b101011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001000010000001  0X0111000X1XXXX01");
    apply_vector ( 24'b111010101001000010000001,17'b0X0111000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101000010000011  111111000X0XXXX00");
    apply_vector ( 24'b010010100101000010000011,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101000010000001  0X0000100X0XXXX00");
    apply_vector ( 24'b111010101101000010000001,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011000010000000  101000100X0XXXX00");
    apply_vector ( 24'b001010100011000010000000,17'b101000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011000010000001  0X0100100X0XXXX00");
    apply_vector ( 24'b111010101011000010000001,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111000010000000  111100100X0XXXX00");
    apply_vector ( 24'b010010100111000010000000,17'b111100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010101111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111000010000000  0X0010100X0XXXX00");
    apply_vector ( 24'b111010101111000010000000,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001100000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000000010000000  100110000X0XXXX00");
    apply_vector ( 24'b001001100000000010000000,17'b100110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000000010000001  0X1110000X1110111");
    apply_vector ( 24'b111001101000000010000001,17'b0X1110000X1110111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100000010000010  110001000X0110110");
    apply_vector ( 24'b010001100100000010000010,17'b110001000X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100000010000000  0X1001000X0110110");
    apply_vector ( 24'b111001101100000010000000,17'b0X1001000X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010000010000001  100101000X0110110");
    apply_vector ( 24'b001001100010000010000001,17'b100101000X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010000010000001  0X1101000X0110110");
    apply_vector ( 24'b111001101010000010000001,17'b0X1101000X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110000010000000  110011000X0110110");
    apply_vector ( 24'b010001100110000010000000,17'b110011000X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110000010000000  0X1011000X0110110");
    apply_vector ( 24'b111001101110000010000000,17'b0X1011000X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001100001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001000010000000  100111000X0110110");
    apply_vector ( 24'b001001100001000010000000,17'b100111000X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001000010000001  0X1111000X1010110");
    apply_vector ( 24'b111001101001000010000001,17'b0X1111000X1010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101000010000011  110000100X0010110");
    apply_vector ( 24'b010001100101000010000011,17'b110000100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101000010000000  0X1000100X0010110");
    apply_vector ( 24'b111001101101000010000000,17'b0X1000100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011000010000001  100100100X0010110");
    apply_vector ( 24'b001001100011000010000001,17'b100100100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011000010000001  0X1100100X0010110");
    apply_vector ( 24'b111001101011000010000001,17'b0X1100100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111000010000000  110010100X0010110");
    apply_vector ( 24'b010001100111000010000000,17'b110010100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111000010000000  0X1010100X0010110");
    apply_vector ( 24'b111001101111000010000000,17'b0X1010100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011100000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000000010000000  101110000X0010110");
    apply_vector ( 24'b001011100000000010000000,17'b101110000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000000010000001  0X0001000X1010111");
    apply_vector ( 24'b111011101000000010000001,17'b0X0001000X1010111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100000010000010  111001000X0010110");
    apply_vector ( 24'b010011100100000010000010,17'b111001000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100000010000001  0X0101000X0010110");
    apply_vector ( 24'b111011101100000010000001,17'b0X0101000X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010000010000001  101101000X0010110");
    apply_vector ( 24'b001011100010000010000001,17'b101101000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010000010000001  0X0011000X0010110");
    apply_vector ( 24'b111011101010000010000001,17'b0X0011000X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110000010000000  111011000X0010110");
    apply_vector ( 24'b010011100110000010000000,17'b111011000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110000010000000  0X0111000X0010110");
    apply_vector ( 24'b111011101110000010000000,17'b0X0111000X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011100001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001000010000000  101111000X0010110");
    apply_vector ( 24'b001011100001000010000000,17'b101111000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001000010000001  0X0000100X1010111");
    apply_vector ( 24'b111011101001000010000001,17'b0X0000100X1010111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101000010000011  111000100X0010110");
    apply_vector ( 24'b010011100101000010000011,17'b111000100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101000010000001  0X0100100X0010110");
    apply_vector ( 24'b111011101101000010000001,17'b0X0100100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011000010000001  101100100X0010110");
    apply_vector ( 24'b001011100011000010000001,17'b101100100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011000010000001  0X0010100X0010110");
    apply_vector ( 24'b111011101011000010000001,17'b0X0010100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111000010000000  111010100X0010110");
    apply_vector ( 24'b010011100111000010000000,17'b111010100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111000010000000  0X0110100X0010110");
    apply_vector ( 24'b111011101111000010000000,17'b0X0110100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000000010000000  100001000X0010110");
    apply_vector ( 24'b001000010000000010000000,17'b100001000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000000010000001  0X1001000X1XXXX01");
    apply_vector ( 24'b111000011000000010000001,17'b0X1001000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100000010000010  110101000X0XXXX00");
    apply_vector ( 24'b010000010100000010000010,17'b110101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100000010000000  0X1101000X0XXXX00");
    apply_vector ( 24'b111000011100000010000000,17'b0X1101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010000010000000  100011000X0XXXX00");
    apply_vector ( 24'b001000010010000010000000,17'b100011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010000010000000  0X1011000X0XXXX00");
    apply_vector ( 24'b111000011010000010000000,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110000010000001  110111000X0XXXX00");
    apply_vector ( 24'b010000010110000010000001,17'b110111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111000011110000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001000010000000  100000100X0XXXX00");
    apply_vector ( 24'b001000010001000010000000,17'b100000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001000010000001  0X1000100X1000111");
    apply_vector ( 24'b111000011001000010000001,17'b0X1000100X1000111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101000010000011  110100100X0000110");
    apply_vector ( 24'b010000010101000010000011,17'b110100100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101000010000000  0X1100100X0000110");
    apply_vector ( 24'b111000011101000010000000,17'b0X1100100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011000010000000  100010100X0000110");
    apply_vector ( 24'b001000010011000010000000,17'b100010100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011000010000000  0X1010100X0000110");
    apply_vector ( 24'b111000011011000010000000,17'b0X1010100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111000010000001  110110100X0000110");
    apply_vector ( 24'b010000010111000010000001,17'b110110100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111000010000000  0X1110100X0000110");
    apply_vector ( 24'b111000011111000010000000,17'b0X1110100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000000010000000  101001000X0000110");
    apply_vector ( 24'b001010010000000010000000,17'b101001000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000000010000001  0X0101000X1XXXX01");
    apply_vector ( 24'b111010011000000010000001,17'b0X0101000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100000010000010  111101000X0XXXX00");
    apply_vector ( 24'b010010010100000010000010,17'b111101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100000010000001  0X0011000X0XXXX00");
    apply_vector ( 24'b111010011100000010000001,17'b0X0011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010000010000000  101011000X0XXXX00");
    apply_vector ( 24'b001010010010000010000000,17'b101011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010000010000000  0X0111000X0XXXX00");
    apply_vector ( 24'b111010011010000010000000,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110000010000001  111111000X0XXXX00");
    apply_vector ( 24'b010010010110000010000001,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110000010000000  0X0000100X0XXXX00");
    apply_vector ( 24'b111010011110000010000000,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001000010000000  101000100X0XXXX00");
    apply_vector ( 24'b001010010001000010000000,17'b101000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001000010000001  0X0100100X1XXXX01");
    apply_vector ( 24'b111010011001000010000001,17'b0X0100100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101000010000011  111100100X0XXXX00");
    apply_vector ( 24'b010010010101000010000011,17'b111100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101000010000001  0X0010100X0XXXX00");
    apply_vector ( 24'b111010011101000010000001,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011000010000000  101010100X0XXXX00");
    apply_vector ( 24'b001010010011000010000000,17'b101010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011000010000000  0X0110100X0XXXX00");
    apply_vector ( 24'b111010011011000010000000,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111000010000001  111110100X0XXXX00");
    apply_vector ( 24'b010010010111000010000001,17'b111110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111000010000000  0X0001100X0XXXX00");
    apply_vector ( 24'b111010011111000010000000,17'b0X0001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000000010000000  100101000X0XXXX00");
    apply_vector ( 24'b001001010000000010000000,17'b100101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000000010000001  0X1101000X1110111");
    apply_vector ( 24'b111001011000000010000001,17'b0X1101000X1110111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100000010000010  110011000X0110110");
    apply_vector ( 24'b010001010100000010000010,17'b110011000X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100000010000000  0X1011000X0110110");
    apply_vector ( 24'b111001011100000010000000,17'b0X1011000X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010000010000001  100111000X0110110");
    apply_vector ( 24'b001001010010000010000001,17'b100111000X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010000010000000  0X1111000X0110110");
    apply_vector ( 24'b111001011010000010000000,17'b0X1111000X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110000010000001  110000100X0110110");
    apply_vector ( 24'b010001010110000010000001,17'b110000100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110000010000000  0X1000100X0110110");
    apply_vector ( 24'b111001011110000010000000,17'b0X1000100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001000010000000  100100100X0110110");
    apply_vector ( 24'b001001010001000010000000,17'b100100100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001000010000001  0X1100100X1XXXX01");
    apply_vector ( 24'b111001011001000010000001,17'b0X1100100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101000010000011  110010100X0XXXX00");
    apply_vector ( 24'b010001010101000010000011,17'b110010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101000010000000  0X1010100X0XXXX00");
    apply_vector ( 24'b111001011101000010000000,17'b0X1010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011000010000001  100110100X0XXXX00");
    apply_vector ( 24'b001001010011000010000001,17'b100110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011000010000000  0X1110100X0XXXX00");
    apply_vector ( 24'b111001011011000010000000,17'b0X1110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111000010000001  110001100X0XXXX00");
    apply_vector ( 24'b010001010111000010000001,17'b110001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111000010000000  0X1001100X0XXXX00");
    apply_vector ( 24'b111001011111000010000000,17'b0X1001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000000010000000  101101000X0XXXX00");
    apply_vector ( 24'b001011010000000010000000,17'b101101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000000010000001  0X0011000X1000011");
    apply_vector ( 24'b111011011000000010000001,17'b0X0011000X1000011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100000010000010  111011000X0000010");
    apply_vector ( 24'b010011010100000010000010,17'b111011000X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100000010000001  0X0111000X0000010");
    apply_vector ( 24'b111011011100000010000001,17'b0X0111000X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010000010000001  101111000X0000010");
    apply_vector ( 24'b001011010010000010000001,17'b101111000X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010000010000000  0X0000100X0000010");
    apply_vector ( 24'b111011011010000010000000,17'b0X0000100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110000010000001  111000100X0000010");
    apply_vector ( 24'b010011010110000010000001,17'b111000100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110000010000000  0X0100100X0000010");
    apply_vector ( 24'b111011011110000010000000,17'b0X0100100X0000010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001000010000000  101100100X0000010");
    apply_vector ( 24'b001011010001000010000000,17'b101100100X0000010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001000010000001  0X0010100X1101111");
    apply_vector ( 24'b111011011001000010000001,17'b0X0010100X1101111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101000010000011  111010100X0101110");
    apply_vector ( 24'b010011010101000010000011,17'b111010100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101000010000001  0X0110100X0101110");
    apply_vector ( 24'b111011011101000010000001,17'b0X0110100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011000010000001  101110100X0101110");
    apply_vector ( 24'b001011010011000010000001,17'b101110100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011000010000000  0X0001100X0101110");
    apply_vector ( 24'b111011011011000010000000,17'b0X0001100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111000010000001  111001100X0101110");
    apply_vector ( 24'b010011010111000010000001,17'b111001100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111000010000000  0X0101100X0101110");
    apply_vector ( 24'b111011011111000010000000,17'b0X0101100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000000010000000  100011000X0101110");
    apply_vector ( 24'b001000110000000010000000,17'b100011000X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000000010000001  0X1011000X1XXXX01");
    apply_vector ( 24'b111000111000000010000001,17'b0X1011000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100000010000010  110111000X0XXXX00");
    apply_vector ( 24'b010000110100000010000010,17'b110111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111000111100000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010000010000000  100000100X0XXXX00");
    apply_vector ( 24'b001000110010000010000000,17'b100000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010000010000001  0X1000100X0XXXX00");
    apply_vector ( 24'b111000111010000010000001,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110000010000001  110100100X0XXXX00");
    apply_vector ( 24'b010000110110000010000001,17'b110100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110000010000000  0X1100100X0XXXX00");
    apply_vector ( 24'b111000111110000010000000,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001000010000000  100010100X0XXXX00");
    apply_vector ( 24'b001000110001000010000000,17'b100010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001000010000001  0X1010100X1XXXX01");
    apply_vector ( 24'b111000111001000010000001,17'b0X1010100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101000010000011  110110100X0XXXX00");
    apply_vector ( 24'b010000110101000010000011,17'b110110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101000010000000  0X1110100X0XXXX00");
    apply_vector ( 24'b111000111101000010000000,17'b0X1110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011000010000000  100001100X0XXXX00");
    apply_vector ( 24'b001000110011000010000000,17'b100001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011000010000001  0X1001100X0XXXX00");
    apply_vector ( 24'b111000111011000010000001,17'b0X1001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111000010000001  110101100X0XXXX00");
    apply_vector ( 24'b010000110111000010000001,17'b110101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111000010000000  0X1101100X0XXXX00");
    apply_vector ( 24'b111000111111000010000000,17'b0X1101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000000010000000  101011000X0XXXX00");
    apply_vector ( 24'b001010110000000010000000,17'b101011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000000010000001  0X0111000X1110111");
    apply_vector ( 24'b111010111000000010000001,17'b0X0111000X1110111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100000010000010  111111000X0110110");
    apply_vector ( 24'b010010110100000010000010,17'b111111000X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100000010000001  0X0000100X0110110");
    apply_vector ( 24'b111010111100000010000001,17'b0X0000100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010000010000000  101000100X0110110");
    apply_vector ( 24'b001010110010000010000000,17'b101000100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010000010000001  0X0100100X0110110");
    apply_vector ( 24'b111010111010000010000001,17'b0X0100100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110000010000001  111100100X0110110");
    apply_vector ( 24'b010010110110000010000001,17'b111100100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110000010000000  0X0010100X0110110");
    apply_vector ( 24'b111010111110000010000000,17'b0X0010100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001000010000000  101010100X0110110");
    apply_vector ( 24'b001010110001000010000000,17'b101010100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001000010000001  0X0110100X1110111");
    apply_vector ( 24'b111010111001000010000001,17'b0X0110100X1110111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101000010000011  111110100X0110110");
    apply_vector ( 24'b010010110101000010000011,17'b111110100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101000010000001  0X0001100X0110110");
    apply_vector ( 24'b111010111101000010000001,17'b0X0001100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011000010000000  101001100X0110110");
    apply_vector ( 24'b001010110011000010000000,17'b101001100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011000010000001  0X0101100X0110110");
    apply_vector ( 24'b111010111011000010000001,17'b0X0101100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111000010000001  111101100X0110110");
    apply_vector ( 24'b010010110111000010000001,17'b111101100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111000010000000  0X0011100X0110110");
    apply_vector ( 24'b111010111111000010000000,17'b0X0011100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000000010000000  100111000X0110110");
    apply_vector ( 24'b001001110000000010000000,17'b100111000X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000000010000001  0X1111000X1110110");
    apply_vector ( 24'b111001111000000010000001,17'b0X1111000X1110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100000010000010  110000100X0110110");
    apply_vector ( 24'b010001110100000010000010,17'b110000100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100000010000000  0X1000100X0110110");
    apply_vector ( 24'b111001111100000010000000,17'b0X1000100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010000010000001  100100100X0110110");
    apply_vector ( 24'b001001110010000010000001,17'b100100100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010000010000001  0X1100100X0110110");
    apply_vector ( 24'b111001111010000010000001,17'b0X1100100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110000010000001  110010100X0110110");
    apply_vector ( 24'b010001110110000010000001,17'b110010100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110000010000000  0X1010100X0110110");
    apply_vector ( 24'b111001111110000010000000,17'b0X1010100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001000010000000  100110100X0110110");
    apply_vector ( 24'b001001110001000010000000,17'b100110100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001000010000001  0X1110100X1010111");
    apply_vector ( 24'b111001111001000010000001,17'b0X1110100X1010111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101000010000011  110001100X0010110");
    apply_vector ( 24'b010001110101000010000011,17'b110001100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101000010000000  0X1001100X0010110");
    apply_vector ( 24'b111001111101000010000000,17'b0X1001100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011000010000001  100101100X0010110");
    apply_vector ( 24'b001001110011000010000001,17'b100101100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011000010000001  0X1101100X0010110");
    apply_vector ( 24'b111001111011000010000001,17'b0X1101100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111000010000001  110011100X0010110");
    apply_vector ( 24'b010001110111000010000001,17'b110011100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111000010000000  0X1011100X0010110");
    apply_vector ( 24'b111001111111000010000000,17'b0X1011100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000000010000000  101111000X0010110");
    apply_vector ( 24'b001011110000000010000000,17'b101111000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000000010000001  0X0000100X1XXXX01");
    apply_vector ( 24'b111011111000000010000001,17'b0X0000100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100000010000010  111000100X0XXXX00");
    apply_vector ( 24'b010011110100000010000010,17'b111000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100000010000001  0X0100100X0XXXX00");
    apply_vector ( 24'b111011111100000010000001,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010000010000001  101100100X0XXXX00");
    apply_vector ( 24'b001011110010000010000001,17'b101100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010000010000001  0X0010100X0XXXX00");
    apply_vector ( 24'b111011111010000010000001,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110000010000001  111010100X0XXXX00");
    apply_vector ( 24'b010011110110000010000001,17'b111010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110000010000000  0X0110100X0XXXX00");
    apply_vector ( 24'b111011111110000010000000,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001000010000000  101110100X0XXXX00");
    apply_vector ( 24'b001011110001000010000000,17'b101110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001000010000001  0X0001100X1XXXX01");
    apply_vector ( 24'b111011111001000010000001,17'b0X0001100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101000010000011  111001100X0XXXX00");
    apply_vector ( 24'b010011110101000010000011,17'b111001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101000010000001  0X0101100X0XXXX00");
    apply_vector ( 24'b111011111101000010000001,17'b0X0101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011000010000001  101101100X0XXXX00");
    apply_vector ( 24'b001011110011000010000001,17'b101101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011000010000001  0X0011100X0XXXX00");
    apply_vector ( 24'b111011111011000010000001,17'b0X0011100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111000010000001  111011100X0XXXX00");
    apply_vector ( 24'b010011110111000010000001,17'b111011100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111000010000000  0X0111100X0XXXX00");
    apply_vector ( 24'b111011111111000010000000,17'b0X0111100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100000000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000000010000000  101000000X0XXXX00");
    apply_vector ( 24'b001100000000000010000000,17'b101000000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000000010000001  0X0100000X1110111");
    apply_vector ( 24'b111100001000000010000001,17'b0X0100000X1110111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100000010000010  111100000X0110110");
    apply_vector ( 24'b010100000100000010000010,17'b111100000X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100000010000000  0X0010000X0110110");
    apply_vector ( 24'b111100001100000010000000,17'b0X0010000X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010000010000000  101010000X0110110");
    apply_vector ( 24'b001100000010000010000000,17'b101010000X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010000010000000  0X0110000X0110110");
    apply_vector ( 24'b111100001010000010000000,17'b0X0110000X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110000010000000  111110000X0110110");
    apply_vector ( 24'b010100000110000010000000,17'b111110000X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110000010000001  0X0001000X0110110");
    apply_vector ( 24'b111100001110000010000001,17'b0X0001000X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001000010000000  101001000X0110110");
    apply_vector ( 24'b001100000001000010000000,17'b101001000X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001000010000001  0X0101000X1001111");
    apply_vector ( 24'b111100001001000010000001,17'b0X0101000X1001111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101000010000011  111101000X0001110");
    apply_vector ( 24'b010100000101000010000011,17'b111101000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101000010000000  0X0011000X0001110");
    apply_vector ( 24'b111100001101000010000000,17'b0X0011000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011000010000000  101011000X0001110");
    apply_vector ( 24'b001100000011000010000000,17'b101011000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011000010000000  0X0111000X0001110");
    apply_vector ( 24'b111100001011000010000000,17'b0X0111000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111000010000000  111111000X0001110");
    apply_vector ( 24'b010100000111000010000000,17'b111111000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111000010000001  0X0000100X0001110");
    apply_vector ( 24'b111100001111000010000001,17'b0X0000100X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110000000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000000010000000  100100000X0001110");
    apply_vector ( 24'b001110000000000010000000,17'b100100000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000000010000001  0X1100000X1001110");
    apply_vector ( 24'b111110001000000010000001,17'b0X1100000X1001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100000010000010  110010000X0001110");
    apply_vector ( 24'b010110000100000010000010,17'b110010000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100000010000001  0X1010000X0001110");
    apply_vector ( 24'b111110001100000010000001,17'b0X1010000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010000010000000  100110000X0001110");
    apply_vector ( 24'b001110000010000010000000,17'b100110000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010000010000000  0X1110000X0001110");
    apply_vector ( 24'b111110001010000010000000,17'b0X1110000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110000010000000  110001000X0001110");
    apply_vector ( 24'b010110000110000010000000,17'b110001000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110000010000001  0X1001000X0001110");
    apply_vector ( 24'b111110001110000010000001,17'b0X1001000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001000010000000  100101000X0001110");
    apply_vector ( 24'b001110000001000010000000,17'b100101000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001000010000001  0X1101000X1XXXX01");
    apply_vector ( 24'b111110001001000010000001,17'b0X1101000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101000010000011  110011000X0XXXX00");
    apply_vector ( 24'b010110000101000010000011,17'b110011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101000010000001  0X1011000X0XXXX00");
    apply_vector ( 24'b111110001101000010000001,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011000010000000  100111000X0XXXX00");
    apply_vector ( 24'b001110000011000010000000,17'b100111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111110001011000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111000010000000  110000100X0XXXX00");
    apply_vector ( 24'b010110000111000010000000,17'b110000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111000010000001  0X1000100X0XXXX00");
    apply_vector ( 24'b111110001111000010000001,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101000000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000000010000000  101100000X0XXXX00");
    apply_vector ( 24'b001101000000000010000000,17'b101100000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000000010000001  0X0010000X1001111");
    apply_vector ( 24'b111101001000000010000001,17'b0X0010000X1001111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100000010000010  111010000X0001110");
    apply_vector ( 24'b010101000100000010000010,17'b111010000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100000010000000  0X0110000X0001110");
    apply_vector ( 24'b111101001100000010000000,17'b0X0110000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010000010000001  101110000X0001110");
    apply_vector ( 24'b001101000010000010000001,17'b101110000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010000010000000  0X0001000X0001110");
    apply_vector ( 24'b111101001010000010000000,17'b0X0001000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110000010000000  111001000X0001110");
    apply_vector ( 24'b010101000110000010000000,17'b111001000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110000010000001  0X0101000X0001110");
    apply_vector ( 24'b111101001110000010000001,17'b0X0101000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001000010000000  101101000X0001110");
    apply_vector ( 24'b001101000001000010000000,17'b101101000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001000010000001  0X0011000X1XXXX01");
    apply_vector ( 24'b111101001001000010000001,17'b0X0011000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101000010000011  111011000X0XXXX00");
    apply_vector ( 24'b010101000101000010000011,17'b111011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101000010000000  0X0111000X0XXXX00");
    apply_vector ( 24'b111101001101000010000000,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011000010000001  101111000X0XXXX00");
    apply_vector ( 24'b001101000011000010000001,17'b101111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011000010000000  0X0000100X0XXXX00");
    apply_vector ( 24'b111101001011000010000000,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111000010000000  111000100X0XXXX00");
    apply_vector ( 24'b010101000111000010000000,17'b111000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111000010000001  0X0100100X0XXXX00");
    apply_vector ( 24'b111101001111000010000001,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111000000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000000010000000  100010000X0XXXX00");
    apply_vector ( 24'b001111000000000010000000,17'b100010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000000010000001  0X1010000X1001111");
    apply_vector ( 24'b111111001000000010000001,17'b0X1010000X1001111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100000010000010  110110000X0001110");
    apply_vector ( 24'b010111000100000010000010,17'b110110000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100000010000001  0X1110000X0001110");
    apply_vector ( 24'b111111001100000010000001,17'b0X1110000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010000010000001  100001000X0001110");
    apply_vector ( 24'b001111000010000010000001,17'b100001000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010000010000000  0X1001000X0001110");
    apply_vector ( 24'b111111001010000010000000,17'b0X1001000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110000010000000  110101000X0001110");
    apply_vector ( 24'b010111000110000010000000,17'b110101000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110000010000001  0X1101000X0001110");
    apply_vector ( 24'b111111001110000010000001,17'b0X1101000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001000010000000  100011000X0001110");
    apply_vector ( 24'b001111000001000010000000,17'b100011000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001000010000001  0X1011000X1101111");
    apply_vector ( 24'b111111001001000010000001,17'b0X1011000X1101111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101000010000011  110111000X0101110");
    apply_vector ( 24'b010111000101000010000011,17'b110111000X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101000010000001  0X1111000X0101110");
    apply_vector ( 24'b111111001101000010000001,17'b0X1111000X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011000010000001  100000100X0101110");
    apply_vector ( 24'b001111000011000010000001,17'b100000100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011000010000000  0X1000100X0101110");
    apply_vector ( 24'b111111001011000010000000,17'b0X1000100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111000010000000  110100100X0101110");
    apply_vector ( 24'b010111000111000010000000,17'b110100100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111000010000001  0X1100100X0101110");
    apply_vector ( 24'b111111001111000010000001,17'b0X1100100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100100000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000000010000000  101010000X0101110");
    apply_vector ( 24'b001100100000000010000000,17'b101010000X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000000010000001  0X0110000X1XXXX01");
    apply_vector ( 24'b111100101000000010000001,17'b0X0110000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100000010000010  111110000X0XXXX00");
    apply_vector ( 24'b010100100100000010000010,17'b111110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100000010000000  0X0001000X0XXXX00");
    apply_vector ( 24'b111100101100000010000000,17'b0X0001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010000010000000  101001000X0XXXX00");
    apply_vector ( 24'b001100100010000010000000,17'b101001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010000010000001  0X0101000X0XXXX00");
    apply_vector ( 24'b111100101010000010000001,17'b0X0101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110000010000000  111101000X0XXXX00");
    apply_vector ( 24'b010100100110000010000000,17'b111101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110000010000001  0X0011000X0XXXX00");
    apply_vector ( 24'b111100101110000010000001,17'b0X0011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100100001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001000010000000  101011000X0XXXX00");
    apply_vector ( 24'b001100100001000010000000,17'b101011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001000010000001  0X0111000X1XXXX01");
    apply_vector ( 24'b111100101001000010000001,17'b0X0111000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101000010000011  111111000X0XXXX00");
    apply_vector ( 24'b010100100101000010000011,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101000010000000  0X0000100X0XXXX00");
    apply_vector ( 24'b111100101101000010000000,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011000010000000  101000100X0XXXX00");
    apply_vector ( 24'b001100100011000010000000,17'b101000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011000010000001  0X0100100X0XXXX00");
    apply_vector ( 24'b111100101011000010000001,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111000010000000  111100100X0XXXX00");
    apply_vector ( 24'b010100100111000010000000,17'b111100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111000010000001  0X0010100X0XXXX00");
    apply_vector ( 24'b111100101111000010000001,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110100000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000000010000000  100110000X0XXXX00");
    apply_vector ( 24'b001110100000000010000000,17'b100110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000000010000001  0X1110000X1001111");
    apply_vector ( 24'b111110101000000010000001,17'b0X1110000X1001111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100000010000010  110001000X0001110");
    apply_vector ( 24'b010110100100000010000010,17'b110001000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100000010000001  0X1001000X0001110");
    apply_vector ( 24'b111110101100000010000001,17'b0X1001000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010000010000000  100101000X0001110");
    apply_vector ( 24'b001110100010000010000000,17'b100101000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010000010000001  0X1101000X0001110");
    apply_vector ( 24'b111110101010000010000001,17'b0X1101000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110000010000000  110011000X0001110");
    apply_vector ( 24'b010110100110000010000000,17'b110011000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110000010000001  0X1011000X0001110");
    apply_vector ( 24'b111110101110000010000001,17'b0X1011000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110100001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001000010000000  100111000X0001110");
    apply_vector ( 24'b001110100001000010000000,17'b100111000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001000010000001  0X1111000X1111111");
    apply_vector ( 24'b111110101001000010000001,17'b0X1111000X1111111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101000010000011  110000100X0111110");
    apply_vector ( 24'b010110100101000010000011,17'b110000100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101000010000001  0X1000100X0111110");
    apply_vector ( 24'b111110101101000010000001,17'b0X1000100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011000010000000  100100100X0111110");
    apply_vector ( 24'b001110100011000010000000,17'b100100100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011000010000001  0X1100100X0111110");
    apply_vector ( 24'b111110101011000010000001,17'b0X1100100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111000010000000  110010100X0111110");
    apply_vector ( 24'b010110100111000010000000,17'b110010100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111000010000001  0X1010100X0111110");
    apply_vector ( 24'b111110101111000010000001,17'b0X1010100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101100000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000000010000000  101110000X0111110");
    apply_vector ( 24'b001101100000000010000000,17'b101110000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000000010000001  0X0001000X1XXXX01");
    apply_vector ( 24'b111101101000000010000001,17'b0X0001000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100000010000010  111001000X0XXXX00");
    apply_vector ( 24'b010101100100000010000010,17'b111001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100000010000000  0X0101000X0XXXX00");
    apply_vector ( 24'b111101101100000010000000,17'b0X0101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010000010000001  101101000X0XXXX00");
    apply_vector ( 24'b001101100010000010000001,17'b101101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010000010000001  0X0011000X0XXXX00");
    apply_vector ( 24'b111101101010000010000001,17'b0X0011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110000010000000  111011000X0XXXX00");
    apply_vector ( 24'b010101100110000010000000,17'b111011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110000010000001  0X0111000X0XXXX00");
    apply_vector ( 24'b111101101110000010000001,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101100001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001000010000000  101111000X0XXXX00");
    apply_vector ( 24'b001101100001000010000000,17'b101111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001000010000001  0X0000100X1010111");
    apply_vector ( 24'b111101101001000010000001,17'b0X0000100X1010111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101000010000011  111000100X0010110");
    apply_vector ( 24'b010101100101000010000011,17'b111000100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101000010000000  0X0100100X0010110");
    apply_vector ( 24'b111101101101000010000000,17'b0X0100100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011000010000001  101100100X0010110");
    apply_vector ( 24'b001101100011000010000001,17'b101100100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011000010000001  0X0010100X0010110");
    apply_vector ( 24'b111101101011000010000001,17'b0X0010100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111000010000000  111010100X0010110");
    apply_vector ( 24'b010101100111000010000000,17'b111010100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111000010000001  0X0110100X0010110");
    apply_vector ( 24'b111101101111000010000001,17'b0X0110100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111100000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000000010000000  100001000X0010110");
    apply_vector ( 24'b001111100000000010000000,17'b100001000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000000010000001  0X1001000X1XXXX01");
    apply_vector ( 24'b111111101000000010000001,17'b0X1001000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100000010000010  110101000X0XXXX00");
    apply_vector ( 24'b010111100100000010000010,17'b110101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100000010000001  0X1101000X0XXXX00");
    apply_vector ( 24'b111111101100000010000001,17'b0X1101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010000010000001  100011000X0XXXX00");
    apply_vector ( 24'b001111100010000010000001,17'b100011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010000010000001  0X1011000X0XXXX00");
    apply_vector ( 24'b111111101010000010000001,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110000010000000  110111000X0XXXX00");
    apply_vector ( 24'b010111100110000010000000,17'b110111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110000010000001  0X1111000X0XXXX00");
    apply_vector ( 24'b111111101110000010000001,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111100001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001000010000000  100000100X0XXXX00");
    apply_vector ( 24'b001111100001000010000000,17'b100000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001000010000001  0X1000100X1XXXX01");
    apply_vector ( 24'b111111101001000010000001,17'b0X1000100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101000010000011  110100100X0XXXX00");
    apply_vector ( 24'b010111100101000010000011,17'b110100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101000010000001  0X1100100X0XXXX00");
    apply_vector ( 24'b111111101101000010000001,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011000010000001  100010100X0XXXX00");
    apply_vector ( 24'b001111100011000010000001,17'b100010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011000010000001  0X1010100X0XXXX00");
    apply_vector ( 24'b111111101011000010000001,17'b0X1010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111000010000000  110110100X0XXXX00");
    apply_vector ( 24'b010111100111000010000000,17'b110110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111000010000001  0X1110100X0XXXX00");
    apply_vector ( 24'b111111101111000010000001,17'b0X1110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000000010000000  101001000X0XXXX00");
    apply_vector ( 24'b001100010000000010000000,17'b101001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000000010000001  0X0101000X1111011");
    apply_vector ( 24'b111100011000000010000001,17'b0X0101000X1111011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100000010000010  111101000X0111010");
    apply_vector ( 24'b010100010100000010000010,17'b111101000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100000010000000  0X0011000X0111010");
    apply_vector ( 24'b111100011100000010000000,17'b0X0011000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010000010000000  101011000X0111010");
    apply_vector ( 24'b001100010010000010000000,17'b101011000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010000010000000  0X0111000X0111010");
    apply_vector ( 24'b111100011010000010000000,17'b0X0111000X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110000010000001  111111000X0111010");
    apply_vector ( 24'b010100010110000010000001,17'b111111000X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110000010000001  0X0000100X0111010");
    apply_vector ( 24'b111100011110000010000001,17'b0X0000100X0111010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001000010000000  101000100X0111010");
    apply_vector ( 24'b001100010001000010000000,17'b101000100X0111010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001000010000001  0X0100100X1XXXX01");
    apply_vector ( 24'b111100011001000010000001,17'b0X0100100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101000010000011  111100100X0XXXX00");
    apply_vector ( 24'b010100010101000010000011,17'b111100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101000010000000  0X0010100X0XXXX00");
    apply_vector ( 24'b111100011101000010000000,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011000010000000  101010100X0XXXX00");
    apply_vector ( 24'b001100010011000010000000,17'b101010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011000010000000  0X0110100X0XXXX00");
    apply_vector ( 24'b111100011011000010000000,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111000010000001  111110100X0XXXX00");
    apply_vector ( 24'b010100010111000010000001,17'b111110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111000010000001  0X0001100X0XXXX00");
    apply_vector ( 24'b111100011111000010000001,17'b0X0001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000000010000000  100101000X0XXXX00");
    apply_vector ( 24'b001110010000000010000000,17'b100101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000000010000001  0X1101000X1001111");
    apply_vector ( 24'b111110011000000010000001,17'b0X1101000X1001111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100000010000010  110011000X0001110");
    apply_vector ( 24'b010110010100000010000010,17'b110011000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100000010000001  0X1011000X0001110");
    apply_vector ( 24'b111110011100000010000001,17'b0X1011000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010000010000000  100111000X0001110");
    apply_vector ( 24'b001110010010000010000000,17'b100111000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010000010000000  0X1111000X0001110");
    apply_vector ( 24'b111110011010000010000000,17'b0X1111000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110000010000001  110000100X0001110");
    apply_vector ( 24'b010110010110000010000001,17'b110000100X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110000010000001  0X1000100X0001110");
    apply_vector ( 24'b111110011110000010000001,17'b0X1000100X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001000010000000  100100100X0001110");
    apply_vector ( 24'b001110010001000010000000,17'b100100100X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001000010000001  0X1100100X1101111");
    apply_vector ( 24'b111110011001000010000001,17'b0X1100100X1101111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101000010000011  110010100X0101110");
    apply_vector ( 24'b010110010101000010000011,17'b110010100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101000010000001  0X1010100X0101110");
    apply_vector ( 24'b111110011101000010000001,17'b0X1010100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011000010000000  100110100X0101110");
    apply_vector ( 24'b001110010011000010000000,17'b100110100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011000010000000  0X1110100X0101110");
    apply_vector ( 24'b111110011011000010000000,17'b0X1110100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111000010000001  110001100X0101110");
    apply_vector ( 24'b010110010111000010000001,17'b110001100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111000010000001  0X1001100X0101110");
    apply_vector ( 24'b111110011111000010000001,17'b0X1001100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000000010000000  101101000X0101110");
    apply_vector ( 24'b001101010000000010000000,17'b101101000X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000000010000001  0X0011000X1XXXX01");
    apply_vector ( 24'b111101011000000010000001,17'b0X0011000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100000010000010  111011000X0XXXX00");
    apply_vector ( 24'b010101010100000010000010,17'b111011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100000010000000  0X0111000X0XXXX00");
    apply_vector ( 24'b111101011100000010000000,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010000010000001  101111000X0XXXX00");
    apply_vector ( 24'b001101010010000010000001,17'b101111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010000010000000  0X0000100X0XXXX00");
    apply_vector ( 24'b111101011010000010000000,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110000010000001  111000100X0XXXX00");
    apply_vector ( 24'b010101010110000010000001,17'b111000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110000010000001  0X0100100X0XXXX00");
    apply_vector ( 24'b111101011110000010000001,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001000010000000  101100100X0XXXX00");
    apply_vector ( 24'b001101010001000010000000,17'b101100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001000010000001  0X0010100X1101111");
    apply_vector ( 24'b111101011001000010000001,17'b0X0010100X1101111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101000010000011  111010100X0101110");
    apply_vector ( 24'b010101010101000010000011,17'b111010100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101000010000000  0X0110100X0101110");
    apply_vector ( 24'b111101011101000010000000,17'b0X0110100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011000010000001  101110100X0101110");
    apply_vector ( 24'b001101010011000010000001,17'b101110100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011000010000000  0X0001100X0101110");
    apply_vector ( 24'b111101011011000010000000,17'b0X0001100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111000010000001  111001100X0101110");
    apply_vector ( 24'b010101010111000010000001,17'b111001100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111000010000001  0X0101100X0101110");
    apply_vector ( 24'b111101011111000010000001,17'b0X0101100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111010000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000000010000000  100011000X0101110");
    apply_vector ( 24'b001111010000000010000000,17'b100011000X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000000010000001  0X1011000X1XXXX01");
    apply_vector ( 24'b111111011000000010000001,17'b0X1011000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100000010000010  110111000X0XXXX00");
    apply_vector ( 24'b010111010100000010000010,17'b110111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100000010000001  0X1111000X0XXXX00");
    apply_vector ( 24'b111111011100000010000001,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010000010000001  100000100X0XXXX00");
    apply_vector ( 24'b001111010010000010000001,17'b100000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010000010000000  0X1000100X0XXXX00");
    apply_vector ( 24'b111111011010000010000000,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110000010000001  110100100X0XXXX00");
    apply_vector ( 24'b010111010110000010000001,17'b110100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110000010000001  0X1100100X0XXXX00");
    apply_vector ( 24'b111111011110000010000001,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111010001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001000010000000  100010100X0XXXX00");
    apply_vector ( 24'b001111010001000010000000,17'b100010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001000010000001  0X1010100X1101110");
    apply_vector ( 24'b111111011001000010000001,17'b0X1010100X1101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101000010000011  110110100X0101110");
    apply_vector ( 24'b010111010101000010000011,17'b110110100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101000010000001  0X1110100X0101110");
    apply_vector ( 24'b111111011101000010000001,17'b0X1110100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011000010000001  100001100X0101110");
    apply_vector ( 24'b001111010011000010000001,17'b100001100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011000010000000  0X1001100X0101110");
    apply_vector ( 24'b111111011011000010000000,17'b0X1001100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111000010000001  110101100X0101110");
    apply_vector ( 24'b010111010111000010000001,17'b110101100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111000010000001  0X1101100X0101110");
    apply_vector ( 24'b111111011111000010000001,17'b0X1101100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000000010000000  101011000X0101110");
    apply_vector ( 24'b001100110000000010000000,17'b101011000X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000000010000001  0X0111000X1101111");
    apply_vector ( 24'b111100111000000010000001,17'b0X0111000X1101111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100000010000010  111111000X0101110");
    apply_vector ( 24'b010100110100000010000010,17'b111111000X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100000010000000  0X0000100X0101110");
    apply_vector ( 24'b111100111100000010000000,17'b0X0000100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010000010000000  101000100X0101110");
    apply_vector ( 24'b001100110010000010000000,17'b101000100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010000010000001  0X0100100X0101110");
    apply_vector ( 24'b111100111010000010000001,17'b0X0100100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110000010000001  111100100X0101110");
    apply_vector ( 24'b010100110110000010000001,17'b111100100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110000010000001  0X0010100X0101110");
    apply_vector ( 24'b111100111110000010000001,17'b0X0010100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001000010000000  101010100X0101110");
    apply_vector ( 24'b001100110001000010000000,17'b101010100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001000010000001  0X0110100X1011011");
    apply_vector ( 24'b111100111001000010000001,17'b0X0110100X1011011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101000010000011  111110100X0011010");
    apply_vector ( 24'b010100110101000010000011,17'b111110100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101000010000000  0X0001100X0011010");
    apply_vector ( 24'b111100111101000010000000,17'b0X0001100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011000010000000  101001100X0011010");
    apply_vector ( 24'b001100110011000010000000,17'b101001100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011000010000001  0X0101100X0011010");
    apply_vector ( 24'b111100111011000010000001,17'b0X0101100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111000010000001  111101100X0011010");
    apply_vector ( 24'b010100110111000010000001,17'b111101100X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111000010000001  0X0011100X0011010");
    apply_vector ( 24'b111100111111000010000001,17'b0X0011100X0011010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000000010000000  100111000X0011010");
    apply_vector ( 24'b001110110000000010000000,17'b100111000X0011010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000000010000001  0X1111000X1XXXX01");
    apply_vector ( 24'b111110111000000010000001,17'b0X1111000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100000010000010  110000100X0XXXX00");
    apply_vector ( 24'b010110110100000010000010,17'b110000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100000010000001  0X1000100X0XXXX00");
    apply_vector ( 24'b111110111100000010000001,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010000010000000  100100100X0XXXX00");
    apply_vector ( 24'b001110110010000010000000,17'b100100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010000010000001  0X1100100X0XXXX00");
    apply_vector ( 24'b111110111010000010000001,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110000010000001  110010100X0XXXX00");
    apply_vector ( 24'b010110110110000010000001,17'b110010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110000010000001  0X1010100X0XXXX00");
    apply_vector ( 24'b111110111110000010000001,17'b0X1010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001000010000000  100110100X0XXXX00");
    apply_vector ( 24'b001110110001000010000000,17'b100110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001000010000001  0X1110100X1XXXX01");
    apply_vector ( 24'b111110111001000010000001,17'b0X1110100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101000010000011  110001100X0XXXX00");
    apply_vector ( 24'b010110110101000010000011,17'b110001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101000010000001  0X1001100X0XXXX00");
    apply_vector ( 24'b111110111101000010000001,17'b0X1001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011000010000000  100101100X0XXXX00");
    apply_vector ( 24'b001110110011000010000000,17'b100101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011000010000001  0X1101100X0XXXX00");
    apply_vector ( 24'b111110111011000010000001,17'b0X1101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111000010000001  110011100X0XXXX00");
    apply_vector ( 24'b010110110111000010000001,17'b110011100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111000010000001  0X1011100X0XXXX00");
    apply_vector ( 24'b111110111111000010000001,17'b0X1011100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000000010000000  101111000X0XXXX00");
    apply_vector ( 24'b001101110000000010000000,17'b101111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000000010000001  0X0000100X1110111");
    apply_vector ( 24'b111101111000000010000001,17'b0X0000100X1110111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100000010000010  111000100X0110110");
    apply_vector ( 24'b010101110100000010000010,17'b111000100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100000010000000  0X0100100X0110110");
    apply_vector ( 24'b111101111100000010000000,17'b0X0100100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010000010000001  101100100X0110110");
    apply_vector ( 24'b001101110010000010000001,17'b101100100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010000010000001  0X0010100X0110110");
    apply_vector ( 24'b111101111010000010000001,17'b0X0010100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110000010000001  111010100X0110110");
    apply_vector ( 24'b010101110110000010000001,17'b111010100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110000010000001  0X0110100X0110110");
    apply_vector ( 24'b111101111110000010000001,17'b0X0110100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001000010000000  101110100X0110110");
    apply_vector ( 24'b001101110001000010000000,17'b101110100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001000010000001  0X0001100X1XXXX01");
    apply_vector ( 24'b111101111001000010000001,17'b0X0001100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101000010000011  111001100X0XXXX00");
    apply_vector ( 24'b010101110101000010000011,17'b111001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101000010000000  0X0101100X0XXXX00");
    apply_vector ( 24'b111101111101000010000000,17'b0X0101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011000010000001  101101100X0XXXX00");
    apply_vector ( 24'b001101110011000010000001,17'b101101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011000010000001  0X0011100X0XXXX00");
    apply_vector ( 24'b111101111011000010000001,17'b0X0011100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111000010000001  111011100X0XXXX00");
    apply_vector ( 24'b010101110111000010000001,17'b111011100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111000010000001  0X0111100X0XXXX00");
    apply_vector ( 24'b111101111111000010000001,17'b0X0111100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111110000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000000010000000  100000100X0XXXX00");
    apply_vector ( 24'b001111110000000010000000,17'b100000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000000010000001  0X1000100X1011111");
    apply_vector ( 24'b111111111000000010000001,17'b0X1000100X1011111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100000010000010  110100100X0011110");
    apply_vector ( 24'b010111110100000010000010,17'b110100100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100000010000001  0X1100100X0011110");
    apply_vector ( 24'b111111111100000010000001,17'b0X1100100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010000010000001  100010100X0011110");
    apply_vector ( 24'b001111110010000010000001,17'b100010100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010000010000001  0X1010100X0011110");
    apply_vector ( 24'b111111111010000010000001,17'b0X1010100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110000010000001  110110100X0011110");
    apply_vector ( 24'b010111110110000010000001,17'b110110100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110000010000001  0X1110100X0011110");
    apply_vector ( 24'b111111111110000010000001,17'b0X1110100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111110001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001000010000000  100001100X0011110");
    apply_vector ( 24'b001111110001000010000000,17'b100001100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001000010000001  0X1001100X1101111");
    apply_vector ( 24'b111111111001000010000001,17'b0X1001100X1101111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101000010000011  110101100X0101110");
    apply_vector ( 24'b010111110101000010000011,17'b110101100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101000010000001  0X1101100X0101110");
    apply_vector ( 24'b111111111101000010000001,17'b0X1101100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011000010000001  100011100X0101110");
    apply_vector ( 24'b001111110011000010000001,17'b100011100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011000010000001  0X1011100X0101110");
    apply_vector ( 24'b111111111011000010000001,17'b0X1011100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111000010000001  110111100X0101110");
    apply_vector ( 24'b010111110111000010000001,17'b110111100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111000010000001  0X1111100X0101110");
    apply_vector ( 24'b111111111111000010000001,17'b0X1111100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000000000000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000000010000000  100000000X0101110");
    apply_vector ( 24'b001000000000000010000000,17'b100000000X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000000010000001  0X1000000X1XXXX01");
    apply_vector ( 24'b111000001000000010000001,17'b0X1000000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100000010000010  110100000X0XXXX00");
    apply_vector ( 24'b010000000100000010000010,17'b110100000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100000010000000  0X1100000X0XXXX00");
    apply_vector ( 24'b111000001100000010000000,17'b0X1100000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010000010000000  100010000X0XXXX00");
    apply_vector ( 24'b001000000010000010000000,17'b100010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010000010000000  0X1010000X0XXXX00");
    apply_vector ( 24'b111000001010000010000000,17'b0X1010000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110000010000000  110110000X0XXXX00");
    apply_vector ( 24'b010000000110000010000000,17'b110110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110000010000000  0X1110000X0XXXX00");
    apply_vector ( 24'b111000001110000010000000,17'b0X1110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001000010000001  100001000X0XXXX00");
    apply_vector ( 24'b001000000001000010000001,17'b100001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001000010000001  0X1001000X1000111");
    apply_vector ( 24'b111000001001000010000001,17'b0X1001000X1000111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101000010000011  110101000X0000110");
    apply_vector ( 24'b010000000101000010000011,17'b110101000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101000010000000  0X1101000X0000110");
    apply_vector ( 24'b111000001101000010000000,17'b0X1101000X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011000010000000  100011000X0000110");
    apply_vector ( 24'b001000000011000010000000,17'b100011000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011000010000000  0X1011000X0000110");
    apply_vector ( 24'b111000001011000010000000,17'b0X1011000X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111000010000000  110111000X0000110");
    apply_vector ( 24'b010000000111000010000000,17'b110111000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000001111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111000010000000  0X1111000X0000110");
    apply_vector ( 24'b111000001111000010000000,17'b0X1111000X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000000010000001  101000000X0000110");
    apply_vector ( 24'b001010000000000010000001,17'b101000000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000000010000001  0X0100000X1XXXX01");
    apply_vector ( 24'b111010001000000010000001,17'b0X0100000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100000010000010  111100000X0XXXX00");
    apply_vector ( 24'b010010000100000010000010,17'b111100000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100000010000001  0X0010000X0XXXX00");
    apply_vector ( 24'b111010001100000010000001,17'b0X0010000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010000010000000  101010000X0XXXX00");
    apply_vector ( 24'b001010000010000010000000,17'b101010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010000010000000  0X0110000X0XXXX00");
    apply_vector ( 24'b111010001010000010000000,17'b0X0110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110000010000000  111110000X0XXXX00");
    apply_vector ( 24'b010010000110000010000000,17'b111110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110000010000000  0X0001000X0XXXX00");
    apply_vector ( 24'b111010001110000010000000,17'b0X0001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001000010000001  101001000X0XXXX00");
    apply_vector ( 24'b001010000001000010000001,17'b101001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001000010000001  0X0101000X1XXXX01");
    apply_vector ( 24'b111010001001000010000001,17'b0X0101000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101000010000011  111101000X0XXXX00");
    apply_vector ( 24'b010010000101000010000011,17'b111101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101000010000001  0X0011000X0XXXX00");
    apply_vector ( 24'b111010001101000010000001,17'b0X0011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011000010000000  101011000X0XXXX00");
    apply_vector ( 24'b001010000011000010000000,17'b101011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011000010000000  0X0111000X0XXXX00");
    apply_vector ( 24'b111010001011000010000000,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111000010000000  111111000X0XXXX00");
    apply_vector ( 24'b010010000111000010000000,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010001111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111000010000000  0X0000100X0XXXX00");
    apply_vector ( 24'b111010001111000010000000,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000000010000001  100100000X0XXXX00");
    apply_vector ( 24'b001001000000000010000001,17'b100100000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000000010000001  0X1100000X1100111");
    apply_vector ( 24'b111001001000000010000001,17'b0X1100000X1100111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100000010000010  110010000X0100110");
    apply_vector ( 24'b010001000100000010000010,17'b110010000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100000010000000  0X1010000X0100110");
    apply_vector ( 24'b111001001100000010000000,17'b0X1010000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010000010000001  100110000X0100110");
    apply_vector ( 24'b001001000010000010000001,17'b100110000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010000010000000  0X1110000X0100110");
    apply_vector ( 24'b111001001010000010000000,17'b0X1110000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110000010000000  110001000X0100110");
    apply_vector ( 24'b010001000110000010000000,17'b110001000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110000010000000  0X1001000X0100110");
    apply_vector ( 24'b111001001110000010000000,17'b0X1001000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001000010000001  100101000X0100110");
    apply_vector ( 24'b001001000001000010000001,17'b100101000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001000010000001  0X1101000X1XXXX01");
    apply_vector ( 24'b111001001001000010000001,17'b0X1101000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101000010000011  110011000X0XXXX00");
    apply_vector ( 24'b010001000101000010000011,17'b110011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101000010000000  0X1011000X0XXXX00");
    apply_vector ( 24'b111001001101000010000000,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011000010000001  100111000X0XXXX00");
    apply_vector ( 24'b001001000011000010000001,17'b100111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111001001011000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111000010000000  110000100X0XXXX00");
    apply_vector ( 24'b010001000111000010000000,17'b110000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001001111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111000010000000  0X1000100X0XXXX00");
    apply_vector ( 24'b111001001111000010000000,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000000010000001  101100000X0XXXX00");
    apply_vector ( 24'b001011000000000010000001,17'b101100000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000000010000001  0X0010000X1100111");
    apply_vector ( 24'b111011001000000010000001,17'b0X0010000X1100111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100000010000010  111010000X0100110");
    apply_vector ( 24'b010011000100000010000010,17'b111010000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100000010000001  0X0110000X0100110");
    apply_vector ( 24'b111011001100000010000001,17'b0X0110000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010000010000001  101110000X0100110");
    apply_vector ( 24'b001011000010000010000001,17'b101110000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010000010000000  0X0001000X0100110");
    apply_vector ( 24'b111011001010000010000000,17'b0X0001000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110000010000000  111001000X0100110");
    apply_vector ( 24'b010011000110000010000000,17'b111001000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110000010000000  0X0101000X0100110");
    apply_vector ( 24'b111011001110000010000000,17'b0X0101000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001000010000001  101101000X0100110");
    apply_vector ( 24'b001011000001000010000001,17'b101101000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001000010000001  0X0011000X1100111");
    apply_vector ( 24'b111011001001000010000001,17'b0X0011000X1100111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101000010000011  111011000X0100110");
    apply_vector ( 24'b010011000101000010000011,17'b111011000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101000010000001  0X0111000X0100110");
    apply_vector ( 24'b111011001101000010000001,17'b0X0111000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011000010000001  101111000X0100110");
    apply_vector ( 24'b001011000011000010000001,17'b101111000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011000010000000  0X0000100X0100110");
    apply_vector ( 24'b111011001011000010000000,17'b0X0000100X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111000010000000  111000100X0100110");
    apply_vector ( 24'b010011000111000010000000,17'b111000100X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011001111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111000010000000  0X0100100X0100110");
    apply_vector ( 24'b111011001111000010000000,17'b0X0100100X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000000010000001  100010000X0100110");
    apply_vector ( 24'b001000100000000010000001,17'b100010000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000000010000001  0X1010000X1100110");
    apply_vector ( 24'b111000101000000010000001,17'b0X1010000X1100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100000010000010  110110000X0100110");
    apply_vector ( 24'b010000100100000010000010,17'b110110000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100000010000000  0X1110000X0100110");
    apply_vector ( 24'b111000101100000010000000,17'b0X1110000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010000010000000  100001000X0100110");
    apply_vector ( 24'b001000100010000010000000,17'b100001000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010000010000001  0X1001000X0100110");
    apply_vector ( 24'b111000101010000010000001,17'b0X1001000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110000010000000  110101000X0100110");
    apply_vector ( 24'b010000100110000010000000,17'b110101000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110000010000000  0X1101000X0100110");
    apply_vector ( 24'b111000101110000010000000,17'b0X1101000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001000010000001  100011000X0100110");
    apply_vector ( 24'b001000100001000010000001,17'b100011000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001000010000001  0X1011000X1XXXX01");
    apply_vector ( 24'b111000101001000010000001,17'b0X1011000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101000010000011  110111000X0XXXX00");
    apply_vector ( 24'b010000100101000010000011,17'b110111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111000101101000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011000010000000  100000100X0XXXX00");
    apply_vector ( 24'b001000100011000010000000,17'b100000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011000010000001  0X1000100X0XXXX00");
    apply_vector ( 24'b111000101011000010000001,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010000100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111000010000000  110100100X0XXXX00");
    apply_vector ( 24'b010000100111000010000000,17'b110100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000101111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111000010000000  0X1100100X0XXXX00");
    apply_vector ( 24'b111000101111000010000000,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000000010000001  101010000X0XXXX00");
    apply_vector ( 24'b001010100000000010000001,17'b101010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000000010000001  0X0110000X1010011");
    apply_vector ( 24'b111010101000000010000001,17'b0X0110000X1010011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100000010000010  111110000X0010010");
    apply_vector ( 24'b010010100100000010000010,17'b111110000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100000010000001  0X0001000X0010010");
    apply_vector ( 24'b111010101100000010000001,17'b0X0001000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010000010000000  101001000X0010010");
    apply_vector ( 24'b001010100010000010000000,17'b101001000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010000010000001  0X0101000X0010010");
    apply_vector ( 24'b111010101010000010000001,17'b0X0101000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110000010000000  111101000X0010010");
    apply_vector ( 24'b010010100110000010000000,17'b111101000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010101110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110000010000000  0X0011000X0010010");
    apply_vector ( 24'b111010101110000010000000,17'b0X0011000X0010010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001000010000001  101011000X0010010");
    apply_vector ( 24'b001010100001000010000001,17'b101011000X0010010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001000010000001  0X0111000X1111111");
    apply_vector ( 24'b111010101001000010000001,17'b0X0111000X1111111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101000010000011  111111000X0111110");
    apply_vector ( 24'b010010100101000010000011,17'b111111000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101000010000001  0X0000100X0111110");
    apply_vector ( 24'b111010101101000010000001,17'b0X0000100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011000010000000  101000100X0111110");
    apply_vector ( 24'b001010100011000010000000,17'b101000100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011000010000001  0X0100100X0111110");
    apply_vector ( 24'b111010101011000010000001,17'b0X0100100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111000010000000  111100100X0111110");
    apply_vector ( 24'b010010100111000010000000,17'b111100100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010101111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111000010000000  0X0010100X0111110");
    apply_vector ( 24'b111010101111000010000000,17'b0X0010100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000000010000001  100110000X0111110");
    apply_vector ( 24'b001001100000000010000001,17'b100110000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000000010000001  0X1110000X1XXXX01");
    apply_vector ( 24'b111001101000000010000001,17'b0X1110000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100000010000010  110001000X0XXXX00");
    apply_vector ( 24'b010001100100000010000010,17'b110001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100000010000000  0X1001000X0XXXX00");
    apply_vector ( 24'b111001101100000010000000,17'b0X1001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010000010000001  100101000X0XXXX00");
    apply_vector ( 24'b001001100010000010000001,17'b100101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010000010000001  0X1101000X0XXXX00");
    apply_vector ( 24'b111001101010000010000001,17'b0X1101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110000010000000  110011000X0XXXX00");
    apply_vector ( 24'b010001100110000010000000,17'b110011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001101110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110000010000000  0X1011000X0XXXX00");
    apply_vector ( 24'b111001101110000010000000,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001000010000001  100111000X0XXXX00");
    apply_vector ( 24'b001001100001000010000001,17'b100111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001000010000001  0X1111000X1010111");
    apply_vector ( 24'b111001101001000010000001,17'b0X1111000X1010111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101000010000011  110000100X0010110");
    apply_vector ( 24'b010001100101000010000011,17'b110000100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101000010000000  0X1000100X0010110");
    apply_vector ( 24'b111001101101000010000000,17'b0X1000100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011000010000001  100100100X0010110");
    apply_vector ( 24'b001001100011000010000001,17'b100100100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011000010000001  0X1100100X0010110");
    apply_vector ( 24'b111001101011000010000001,17'b0X1100100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111000010000000  110010100X0010110");
    apply_vector ( 24'b010001100111000010000000,17'b110010100X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001101111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111000010000000  0X1010100X0010110");
    apply_vector ( 24'b111001101111000010000000,17'b0X1010100X0010110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000000010000001  101110000X0010110");
    apply_vector ( 24'b001011100000000010000001,17'b101110000X0010110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000000010000001  0X0001000X1XXXX01");
    apply_vector ( 24'b111011101000000010000001,17'b0X0001000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100000010000010  111001000X0XXXX00");
    apply_vector ( 24'b010011100100000010000010,17'b111001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100000010000001  0X0101000X0XXXX00");
    apply_vector ( 24'b111011101100000010000001,17'b0X0101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010000010000001  101101000X0XXXX00");
    apply_vector ( 24'b001011100010000010000001,17'b101101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010000010000001  0X0011000X0XXXX00");
    apply_vector ( 24'b111011101010000010000001,17'b0X0011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110000010000000  111011000X0XXXX00");
    apply_vector ( 24'b010011100110000010000000,17'b111011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011101110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110000010000000  0X0111000X0XXXX00");
    apply_vector ( 24'b111011101110000010000000,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001000010000001  101111000X0XXXX00");
    apply_vector ( 24'b001011100001000010000001,17'b101111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001000010000001  0X0000100X1XXXX01");
    apply_vector ( 24'b111011101001000010000001,17'b0X0000100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101000010000011  111000100X0XXXX00");
    apply_vector ( 24'b010011100101000010000011,17'b111000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101000010000001  0X0100100X0XXXX00");
    apply_vector ( 24'b111011101101000010000001,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011000010000001  101100100X0XXXX00");
    apply_vector ( 24'b001011100011000010000001,17'b101100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011000010000001  0X0010100X0XXXX00");
    apply_vector ( 24'b111011101011000010000001,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111000010000000  111010100X0XXXX00");
    apply_vector ( 24'b010011100111000010000000,17'b111010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011101111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111000010000000  0X0110100X0XXXX00");
    apply_vector ( 24'b111011101111000010000000,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000000010000001  100001000X0XXXX00");
    apply_vector ( 24'b001000010000000010000001,17'b100001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000000010000001  0X1001000X1100111");
    apply_vector ( 24'b111000011000000010000001,17'b0X1001000X1100111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100000010000010  110101000X0100110");
    apply_vector ( 24'b010000010100000010000010,17'b110101000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100000010000000  0X1101000X0100110");
    apply_vector ( 24'b111000011100000010000000,17'b0X1101000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010000010000000  100011000X0100110");
    apply_vector ( 24'b001000010010000010000000,17'b100011000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010000010000000  0X1011000X0100110");
    apply_vector ( 24'b111000011010000010000000,17'b0X1011000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110000010000001  110111000X0100110");
    apply_vector ( 24'b010000010110000010000001,17'b110111000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110000010000000  0X1111000X0100110");
    apply_vector ( 24'b111000011110000010000000,17'b0X1111000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001000010000001  100000100X0100110");
    apply_vector ( 24'b001000010001000010000001,17'b100000100X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001000010000001  0X1000100X1000110");
    apply_vector ( 24'b111000011001000010000001,17'b0X1000100X1000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101000010000011  110100100X0000110");
    apply_vector ( 24'b010000010101000010000011,17'b110100100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101000010000000  0X1100100X0000110");
    apply_vector ( 24'b111000011101000010000000,17'b0X1100100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011000010000000  100010100X0000110");
    apply_vector ( 24'b001000010011000010000000,17'b100010100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011000010000000  0X1010100X0000110");
    apply_vector ( 24'b111000011011000010000000,17'b0X1010100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111000010000001  110110100X0000110");
    apply_vector ( 24'b010000010111000010000001,17'b110110100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111000010000000  0X1110100X0000110");
    apply_vector ( 24'b111000011111000010000000,17'b0X1110100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000000010000001  101001000X0000110");
    apply_vector ( 24'b001010010000000010000001,17'b101001000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000000010000001  0X0101000X1000111");
    apply_vector ( 24'b111010011000000010000001,17'b0X0101000X1000111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100000010000010  111101000X0000110");
    apply_vector ( 24'b010010010100000010000010,17'b111101000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100000010000001  0X0011000X0000110");
    apply_vector ( 24'b111010011100000010000001,17'b0X0011000X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010000010000000  101011000X0000110");
    apply_vector ( 24'b001010010010000010000000,17'b101011000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010000010000000  0X0111000X0000110");
    apply_vector ( 24'b111010011010000010000000,17'b0X0111000X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110000010000001  111111000X0000110");
    apply_vector ( 24'b010010010110000010000001,17'b111111000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110000010000000  0X0000100X0000110");
    apply_vector ( 24'b111010011110000010000000,17'b0X0000100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001000010000001  101000100X0000110");
    apply_vector ( 24'b001010010001000010000001,17'b101000100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001000010000001  0X0100100X1000111");
    apply_vector ( 24'b111010011001000010000001,17'b0X0100100X1000111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101000010000011  111100100X0000110");
    apply_vector ( 24'b010010010101000010000011,17'b111100100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101000010000001  0X0010100X0000110");
    apply_vector ( 24'b111010011101000010000001,17'b0X0010100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011000010000000  101010100X0000110");
    apply_vector ( 24'b001010010011000010000000,17'b101010100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011000010000000  0X0110100X0000110");
    apply_vector ( 24'b111010011011000010000000,17'b0X0110100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010010010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111000010000001  111110100X0000110");
    apply_vector ( 24'b010010010111000010000001,17'b111110100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111000010000000  0X0001100X0000110");
    apply_vector ( 24'b111010011111000010000000,17'b0X0001100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000000010000001  100101000X0000110");
    apply_vector ( 24'b001001010000000010000001,17'b100101000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000000010000001  0X1101000X1XXXX01");
    apply_vector ( 24'b111001011000000010000001,17'b0X1101000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100000010000010  110011000X0XXXX00");
    apply_vector ( 24'b010001010100000010000010,17'b110011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100000010000000  0X1011000X0XXXX00");
    apply_vector ( 24'b111001011100000010000000,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010000010000001  100111000X0XXXX00");
    apply_vector ( 24'b001001010010000010000001,17'b100111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111001011010000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110000010000001  110000100X0XXXX00");
    apply_vector ( 24'b010001010110000010000001,17'b110000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110000010000000  0X1000100X0XXXX00");
    apply_vector ( 24'b111001011110000010000000,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001000010000001  100100100X0XXXX00");
    apply_vector ( 24'b001001010001000010000001,17'b100100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001000010000001  0X1100100X1000111");
    apply_vector ( 24'b111001011001000010000001,17'b0X1100100X1000111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101000010000011  110010100X0000110");
    apply_vector ( 24'b010001010101000010000011,17'b110010100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101000010000000  0X1010100X0000110");
    apply_vector ( 24'b111001011101000010000000,17'b0X1010100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011000010000001  100110100X0000110");
    apply_vector ( 24'b001001010011000010000001,17'b100110100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011000010000000  0X1110100X0000110");
    apply_vector ( 24'b111001011011000010000000,17'b0X1110100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111000010000001  110001100X0000110");
    apply_vector ( 24'b010001010111000010000001,17'b110001100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111000010000000  0X1001100X0000110");
    apply_vector ( 24'b111001011111000010000000,17'b0X1001100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000000010000001  101101000X0000110");
    apply_vector ( 24'b001011010000000010000001,17'b101101000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000000010000001  0X0011000X1XXXX01");
    apply_vector ( 24'b111011011000000010000001,17'b0X0011000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100000010000010  111011000X0XXXX00");
    apply_vector ( 24'b010011010100000010000010,17'b111011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100000010000001  0X0111000X0XXXX00");
    apply_vector ( 24'b111011011100000010000001,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010000010000001  101111000X0XXXX00");
    apply_vector ( 24'b001011010010000010000001,17'b101111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010000010000000  0X0000100X0XXXX00");
    apply_vector ( 24'b111011011010000010000000,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110000010000001  111000100X0XXXX00");
    apply_vector ( 24'b010011010110000010000001,17'b111000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011011110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110000010000000  0X0100100X0XXXX00");
    apply_vector ( 24'b111011011110000010000000,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001000010000001  101100100X0XXXX00");
    apply_vector ( 24'b001011010001000010000001,17'b101100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001000010000001  0X0010100X1XXXX01");
    apply_vector ( 24'b111011011001000010000001,17'b0X0010100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101000010000011  111010100X0XXXX00");
    apply_vector ( 24'b010011010101000010000011,17'b111010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101000010000001  0X0110100X0XXXX00");
    apply_vector ( 24'b111011011101000010000001,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011000010000001  101110100X0XXXX00");
    apply_vector ( 24'b001011010011000010000001,17'b101110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011000010000000  0X0001100X0XXXX00");
    apply_vector ( 24'b111011011011000010000000,17'b0X0001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010011010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111000010000001  111001100X0XXXX00");
    apply_vector ( 24'b010011010111000010000001,17'b111001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011011111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111000010000000  0X0101100X0XXXX00");
    apply_vector ( 24'b111011011111000010000000,17'b0X0101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000000010000001  100011000X0XXXX00");
    apply_vector ( 24'b001000110000000010000001,17'b100011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000000010000001  0X1011000X1100111");
    apply_vector ( 24'b111000111000000010000001,17'b0X1011000X1100111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100000010000010  110111000X0100110");
    apply_vector ( 24'b010000110100000010000010,17'b110111000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100000010000000  0X1111000X0100110");
    apply_vector ( 24'b111000111100000010000000,17'b0X1111000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010000010000000  100000100X0100110");
    apply_vector ( 24'b001000110010000010000000,17'b100000100X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010000010000001  0X1000100X0100110");
    apply_vector ( 24'b111000111010000010000001,17'b0X1000100X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110000010000001  110100100X0100110");
    apply_vector ( 24'b010000110110000010000001,17'b110100100X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110000010000000  0X1100100X0100110");
    apply_vector ( 24'b111000111110000010000000,17'b0X1100100X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001000010000001  100010100X0100110");
    apply_vector ( 24'b001000110001000010000001,17'b100010100X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001000010000001  0X1010100X1000111");
    apply_vector ( 24'b111000111001000010000001,17'b0X1010100X1000111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101000010000011  110110100X0000110");
    apply_vector ( 24'b010000110101000010000011,17'b110110100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101000010000000  0X1110100X0000110");
    apply_vector ( 24'b111000111101000010000000,17'b0X1110100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011000010000000  100001100X0000110");
    apply_vector ( 24'b001000110011000010000000,17'b100001100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011000010000001  0X1001100X0000110");
    apply_vector ( 24'b111000111011000010000001,17'b0X1001100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111000010000001  110101100X0000110");
    apply_vector ( 24'b010000110111000010000001,17'b110101100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111000010000000  0X1101100X0000110");
    apply_vector ( 24'b111000111111000010000000,17'b0X1101100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001010110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000000010000001  101011000X0000110");
    apply_vector ( 24'b001010110000000010000001,17'b101011000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111010111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000000010000001  0X0111000X1XXXX01");
    apply_vector ( 24'b111010111000000010000001,17'b0X0111000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100000010000010  111111000X0XXXX00");
    apply_vector ( 24'b010010110100000010000010,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100000010000001  0X0000100X0XXXX00");
    apply_vector ( 24'b111010111100000010000001,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010000010000000  101000100X0XXXX00");
    apply_vector ( 24'b001010110010000010000000,17'b101000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010000010000001  0X0100100X0XXXX00");
    apply_vector ( 24'b111010111010000010000001,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110000010000001  111100100X0XXXX00");
    apply_vector ( 24'b010010110110000010000001,17'b111100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110000010000000  0X0010100X0XXXX00");
    apply_vector ( 24'b111010111110000010000000,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001000010000001  101010100X0XXXX00");
    apply_vector ( 24'b001010110001000010000001,17'b101010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001000010000001  0X0110100X1XXXX01");
    apply_vector ( 24'b111010111001000010000001,17'b0X0110100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101000010000011  111110100X0XXXX00");
    apply_vector ( 24'b010010110101000010000011,17'b111110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101000010000001  0X0001100X0XXXX00");
    apply_vector ( 24'b111010111101000010000001,17'b0X0001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001010110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011000010000000  101001100X0XXXX00");
    apply_vector ( 24'b001010110011000010000000,17'b101001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011000010000001  0X0101100X0XXXX00");
    apply_vector ( 24'b111010111011000010000001,17'b0X0101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010010110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111000010000001  111101100X0XXXX00");
    apply_vector ( 24'b010010110111000010000001,17'b111101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111010111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111000010000000  0X0011100X0XXXX00");
    apply_vector ( 24'b111010111111000010000000,17'b0X0011100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000000010000001  100111000X0XXXX00");
    apply_vector ( 24'b001001110000000010000001,17'b100111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000000010000001  0X1111000X1110111");
    apply_vector ( 24'b111001111000000010000001,17'b0X1111000X1110111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100000010000010  110000100X0110110");
    apply_vector ( 24'b010001110100000010000010,17'b110000100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100000010000000  0X1000100X0110110");
    apply_vector ( 24'b111001111100000010000000,17'b0X1000100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010000010000001  100100100X0110110");
    apply_vector ( 24'b001001110010000010000001,17'b100100100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010000010000001  0X1100100X0110110");
    apply_vector ( 24'b111001111010000010000001,17'b0X1100100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010001110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110000010000001  110010100X0110110");
    apply_vector ( 24'b010001110110000010000001,17'b110010100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110000010000000  0X1010100X0110110");
    apply_vector ( 24'b111001111110000010000000,17'b0X1010100X0110110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001001110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001000010000001  100110100X0110110");
    apply_vector ( 24'b001001110001000010000001,17'b100110100X0110110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111001111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001000010000001  0X1110100X1XXXX01");
    apply_vector ( 24'b111001111001000010000001,17'b0X1110100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101000010000011  110001100X0XXXX00");
    apply_vector ( 24'b010001110101000010000011,17'b110001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101000010000000  0X1001100X0XXXX00");
    apply_vector ( 24'b111001111101000010000000,17'b0X1001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001001110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011000010000001  100101100X0XXXX00");
    apply_vector ( 24'b001001110011000010000001,17'b100101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011000010000001  0X1101100X0XXXX00");
    apply_vector ( 24'b111001111011000010000001,17'b0X1101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010001110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111000010000001  110011100X0XXXX00");
    apply_vector ( 24'b010001110111000010000001,17'b110011100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111001111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111000010000000  0X1011100X0XXXX00");
    apply_vector ( 24'b111001111111000010000000,17'b0X1011100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001011110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000000010000001  101111000X0XXXX00");
    apply_vector ( 24'b001011110000000010000001,17'b101111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111011111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000000010000001  0X0000100X1011111");
    apply_vector ( 24'b111011111000000010000001,17'b0X0000100X1011111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100000010000010  111000100X0011110");
    apply_vector ( 24'b010011110100000010000010,17'b111000100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100000010000001  0X0100100X0011110");
    apply_vector ( 24'b111011111100000010000001,17'b0X0100100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010000010000001  101100100X0011110");
    apply_vector ( 24'b001011110010000010000001,17'b101100100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010000010000001  0X0010100X0011110");
    apply_vector ( 24'b111011111010000010000001,17'b0X0010100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110000010000001  111010100X0011110");
    apply_vector ( 24'b010011110110000010000001,17'b111010100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110000010000000  0X0110100X0011110");
    apply_vector ( 24'b111011111110000010000000,17'b0X0110100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001000010000001  101110100X0011110");
    apply_vector ( 24'b001011110001000010000001,17'b101110100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001000010000001  0X0001100X1110011");
    apply_vector ( 24'b111011111001000010000001,17'b0X0001100X1110011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101000010000011  111001100X0110010");
    apply_vector ( 24'b010011110101000010000011,17'b111001100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101000010000001  0X0101100X0110010");
    apply_vector ( 24'b111011111101000010000001,17'b0X0101100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001011110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011000010000001  101101100X0110010");
    apply_vector ( 24'b001011110011000010000001,17'b101101100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011000010000001  0X0011100X0110010");
    apply_vector ( 24'b111011111011000010000001,17'b0X0011100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010011110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111000010000001  111011100X0110010");
    apply_vector ( 24'b010011110111000010000001,17'b111011100X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111011111111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111000010000000  0X0111100X0110010");
    apply_vector ( 24'b111011111111000010000000,17'b0X0111100X0110010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000000010000001  101000000X0110010");
    apply_vector ( 24'b001100000000000010000001,17'b101000000X0110010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000000010000001  0X0100000X1XXXX01");
    apply_vector ( 24'b111100001000000010000001,17'b0X0100000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100000010000010  111100000X0XXXX00");
    apply_vector ( 24'b010100000100000010000010,17'b111100000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100000010000000  0X0010000X0XXXX00");
    apply_vector ( 24'b111100001100000010000000,17'b0X0010000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010000010000000  101010000X0XXXX00");
    apply_vector ( 24'b001100000010000010000000,17'b101010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010000010000000  0X0110000X0XXXX00");
    apply_vector ( 24'b111100001010000010000000,17'b0X0110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110000010000000  111110000X0XXXX00");
    apply_vector ( 24'b010100000110000010000000,17'b111110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110000010000001  0X0001000X0XXXX00");
    apply_vector ( 24'b111100001110000010000001,17'b0X0001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001000010000001  101001000X0XXXX00");
    apply_vector ( 24'b001100000001000010000001,17'b101001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001000010000001  0X0101000X1XXXX01");
    apply_vector ( 24'b111100001001000010000001,17'b0X0101000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101000010000011  111101000X0XXXX00");
    apply_vector ( 24'b010100000101000010000011,17'b111101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101000010000000  0X0011000X0XXXX00");
    apply_vector ( 24'b111100001101000010000000,17'b0X0011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011000010000000  101011000X0XXXX00");
    apply_vector ( 24'b001100000011000010000000,17'b101011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011000010000000  0X0111000X0XXXX00");
    apply_vector ( 24'b111100001011000010000000,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111000010000000  111111000X0XXXX00");
    apply_vector ( 24'b010100000111000010000000,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111000010000001  0X0000100X0XXXX00");
    apply_vector ( 24'b111100001111000010000001,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000000010000001  100100000X0XXXX00");
    apply_vector ( 24'b001110000000000010000001,17'b100100000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000000010000001  0X1100000X1001111");
    apply_vector ( 24'b111110001000000010000001,17'b0X1100000X1001111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100000010000010  110010000X0001110");
    apply_vector ( 24'b010110000100000010000010,17'b110010000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100000010000001  0X1010000X0001110");
    apply_vector ( 24'b111110001100000010000001,17'b0X1010000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010000010000000  100110000X0001110");
    apply_vector ( 24'b001110000010000010000000,17'b100110000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010000010000000  0X1110000X0001110");
    apply_vector ( 24'b111110001010000010000000,17'b0X1110000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110000010000000  110001000X0001110");
    apply_vector ( 24'b010110000110000010000000,17'b110001000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110000010000001  0X1001000X0001110");
    apply_vector ( 24'b111110001110000010000001,17'b0X1001000X0001110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001000010000001  100101000X0001110");
    apply_vector ( 24'b001110000001000010000001,17'b100101000X0001110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001000010000001  0X1101000X1111111");
    apply_vector ( 24'b111110001001000010000001,17'b0X1101000X1111111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101000010000011  110011000X0111110");
    apply_vector ( 24'b010110000101000010000011,17'b110011000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101000010000001  0X1011000X0111110");
    apply_vector ( 24'b111110001101000010000001,17'b0X1011000X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110000011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011000010000000  100111000X0111110");
    apply_vector ( 24'b001110000011000010000000,17'b100111000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011000010000000  0X1111000X0111110");
    apply_vector ( 24'b111110001011000010000000,17'b0X1111000X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111000010000000  110000100X0111110");
    apply_vector ( 24'b010110000111000010000000,17'b110000100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111000010000001  0X1000100X0111110");
    apply_vector ( 24'b111110001111000010000001,17'b0X1000100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000000010000001  101100000X0111110");
    apply_vector ( 24'b001101000000000010000001,17'b101100000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000000010000001  0X0010000X1XXXX01");
    apply_vector ( 24'b111101001000000010000001,17'b0X0010000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100000010000010  111010000X0XXXX00");
    apply_vector ( 24'b010101000100000010000010,17'b111010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100000010000000  0X0110000X0XXXX00");
    apply_vector ( 24'b111101001100000010000000,17'b0X0110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010000010000001  101110000X0XXXX00");
    apply_vector ( 24'b001101000010000010000001,17'b101110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010000010000000  0X0001000X0XXXX00");
    apply_vector ( 24'b111101001010000010000000,17'b0X0001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110000010000000  111001000X0XXXX00");
    apply_vector ( 24'b010101000110000010000000,17'b111001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110000010000001  0X0101000X0XXXX00");
    apply_vector ( 24'b111101001110000010000001,17'b0X0101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001000010000001  101101000X0XXXX00");
    apply_vector ( 24'b001101000001000010000001,17'b101101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001000010000001  0X0011000X1001011");
    apply_vector ( 24'b111101001001000010000001,17'b0X0011000X1001011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101000010000011  111011000X0001010");
    apply_vector ( 24'b010101000101000010000011,17'b111011000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101000010000000  0X0111000X0001010");
    apply_vector ( 24'b111101001101000010000000,17'b0X0111000X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011000010000001  101111000X0001010");
    apply_vector ( 24'b001101000011000010000001,17'b101111000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011000010000000  0X0000100X0001010");
    apply_vector ( 24'b111101001011000010000000,17'b0X0000100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111000010000000  111000100X0001010");
    apply_vector ( 24'b010101000111000010000000,17'b111000100X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111000010000001  0X0100100X0001010");
    apply_vector ( 24'b111101001111000010000001,17'b0X0100100X0001010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000000010000001  100010000X0001010");
    apply_vector ( 24'b001111000000000010000001,17'b100010000X0001010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000000010000001  0X1010000X1XXXX01");
    apply_vector ( 24'b111111001000000010000001,17'b0X1010000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111000100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100000010000010  110110000X0XXXX00");
    apply_vector ( 24'b010111000100000010000010,17'b110110000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100000010000001  0X1110000X0XXXX00");
    apply_vector ( 24'b111111001100000010000001,17'b0X1110000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111000010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010000010000001  100001000X0XXXX00");
    apply_vector ( 24'b001111000010000010000001,17'b100001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010000010000000  0X1001000X0XXXX00");
    apply_vector ( 24'b111111001010000010000000,17'b0X1001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110000010000000  110101000X0XXXX00");
    apply_vector ( 24'b010111000110000010000000,17'b110101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110000010000001  0X1101000X0XXXX00");
    apply_vector ( 24'b111111001110000010000001,17'b0X1101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111000001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001000010000001  100011000X0XXXX00");
    apply_vector ( 24'b001111000001000010000001,17'b100011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001000010000001  0X1011000X1XXXX01");
    apply_vector ( 24'b111111001001000010000001,17'b0X1011000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111000101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101000010000011  110111000X0XXXX00");
    apply_vector ( 24'b010111000101000010000011,17'b110111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101000010000001  0X1111000X0XXXX00");
    apply_vector ( 24'b111111001101000010000001,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111000011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011000010000001  100000100X0XXXX00");
    apply_vector ( 24'b001111000011000010000001,17'b100000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011000010000000  0X1000100X0XXXX00");
    apply_vector ( 24'b111111001011000010000000,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111000111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111000010000000  110100100X0XXXX00");
    apply_vector ( 24'b010111000111000010000000,17'b110100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111001111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111000010000001  0X1100100X0XXXX00");
    apply_vector ( 24'b111111001111000010000001,17'b0X1100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000000010000001  101010000X0XXXX00");
    apply_vector ( 24'b001100100000000010000001,17'b101010000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000000010000001  0X0110000X1100111");
    apply_vector ( 24'b111100101000000010000001,17'b0X0110000X1100111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100000010000010  111110000X0100110");
    apply_vector ( 24'b010100100100000010000010,17'b111110000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100000010000000  0X0001000X0100110");
    apply_vector ( 24'b111100101100000010000000,17'b0X0001000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010000010000000  101001000X0100110");
    apply_vector ( 24'b001100100010000010000000,17'b101001000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010000010000001  0X0101000X0100110");
    apply_vector ( 24'b111100101010000010000001,17'b0X0101000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110000010000000  111101000X0100110");
    apply_vector ( 24'b010100100110000010000000,17'b111101000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110000010000001  0X0011000X0100110");
    apply_vector ( 24'b111100101110000010000001,17'b0X0011000X0100110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001000010000001  101011000X0100110");
    apply_vector ( 24'b001100100001000010000001,17'b101011000X0100110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001000010000001  0X0111000X1111111");
    apply_vector ( 24'b111100101001000010000001,17'b0X0111000X1111111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101000010000011  111111000X0111110");
    apply_vector ( 24'b010100100101000010000011,17'b111111000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101000010000000  0X0000100X0111110");
    apply_vector ( 24'b111100101101000010000000,17'b0X0000100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011000010000000  101000100X0111110");
    apply_vector ( 24'b001100100011000010000000,17'b101000100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011000010000001  0X0100100X0111110");
    apply_vector ( 24'b111100101011000010000001,17'b0X0100100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111000010000000  111100100X0111110");
    apply_vector ( 24'b010100100111000010000000,17'b111100100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111000010000001  0X0010100X0111110");
    apply_vector ( 24'b111100101111000010000001,17'b0X0010100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000000010000001  100110000X0111110");
    apply_vector ( 24'b001110100000000010000001,17'b100110000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000000010000001  0X1110000X1XXXX01");
    apply_vector ( 24'b111110101000000010000001,17'b0X1110000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100000010000010  110001000X0XXXX00");
    apply_vector ( 24'b010110100100000010000010,17'b110001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100000010000001  0X1001000X0XXXX00");
    apply_vector ( 24'b111110101100000010000001,17'b0X1001000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110100010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010000010000000  100101000X0XXXX00");
    apply_vector ( 24'b001110100010000010000000,17'b100101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010000010000001  0X1101000X0XXXX00");
    apply_vector ( 24'b111110101010000010000001,17'b0X1101000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110000010000000  110011000X0XXXX00");
    apply_vector ( 24'b010110100110000010000000,17'b110011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110000010000001  0X1011000X0XXXX00");
    apply_vector ( 24'b111110101110000010000001,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001000010000001  100111000X0XXXX00");
    apply_vector ( 24'b001110100001000010000001,17'b100111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001000010000001  0X1111000X1111110");
    apply_vector ( 24'b111110101001000010000001,17'b0X1111000X1111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101000010000011  110000100X0111110");
    apply_vector ( 24'b010110100101000010000011,17'b110000100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101000010000001  0X1000100X0111110");
    apply_vector ( 24'b111110101101000010000001,17'b0X1000100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110100011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011000010000000  100100100X0111110");
    apply_vector ( 24'b001110100011000010000000,17'b100100100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011000010000001  0X1100100X0111110");
    apply_vector ( 24'b111110101011000010000001,17'b0X1100100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111000010000000  110010100X0111110");
    apply_vector ( 24'b010110100111000010000000,17'b110010100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111000010000001  0X1010100X0111110");
    apply_vector ( 24'b111110101111000010000001,17'b0X1010100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000000010000001  101110000X0111110");
    apply_vector ( 24'b001101100000000010000001,17'b101110000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000000010000001  0X0001000X1111111");
    apply_vector ( 24'b111101101000000010000001,17'b0X0001000X1111111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100000010000010  111001000X0111110");
    apply_vector ( 24'b010101100100000010000010,17'b111001000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100000010000000  0X0101000X0111110");
    apply_vector ( 24'b111101101100000010000000,17'b0X0101000X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010000010000001  101101000X0111110");
    apply_vector ( 24'b001101100010000010000001,17'b101101000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010000010000001  0X0011000X0111110");
    apply_vector ( 24'b111101101010000010000001,17'b0X0011000X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110000010000000  111011000X0111110");
    apply_vector ( 24'b010101100110000010000000,17'b111011000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110000010000001  0X0111000X0111110");
    apply_vector ( 24'b111101101110000010000001,17'b0X0111000X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001000010000001  101111000X0111110");
    apply_vector ( 24'b001101100001000010000001,17'b101111000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001000010000001  0X0000100X1XXXX01");
    apply_vector ( 24'b111101101001000010000001,17'b0X0000100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101000010000011  111000100X0XXXX00");
    apply_vector ( 24'b010101100101000010000011,17'b111000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101000010000000  0X0100100X0XXXX00");
    apply_vector ( 24'b111101101101000010000000,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011000010000001  101100100X0XXXX00");
    apply_vector ( 24'b001101100011000010000001,17'b101100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011000010000001  0X0010100X0XXXX00");
    apply_vector ( 24'b111101101011000010000001,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111000010000000  111010100X0XXXX00");
    apply_vector ( 24'b010101100111000010000000,17'b111010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111000010000001  0X0110100X0XXXX00");
    apply_vector ( 24'b111101101111000010000001,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111100000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000000010000001  100001000X0XXXX00");
    apply_vector ( 24'b001111100000000010000001,17'b100001000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111101000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000000010000001  0X1001000X1011111");
    apply_vector ( 24'b111111101000000010000001,17'b0X1001000X1011111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111100100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100000010000010  110101000X0011110");
    apply_vector ( 24'b010111100100000010000010,17'b110101000X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100000010000001  0X1101000X0011110");
    apply_vector ( 24'b111111101100000010000001,17'b0X1101000X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111100010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010000010000001  100011000X0011110");
    apply_vector ( 24'b001111100010000010000001,17'b100011000X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010000010000001  0X1011000X0011110");
    apply_vector ( 24'b111111101010000010000001,17'b0X1011000X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111100110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110000010000000  110111000X0011110");
    apply_vector ( 24'b010111100110000010000000,17'b110111000X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110000010000001  0X1111000X0011110");
    apply_vector ( 24'b111111101110000010000001,17'b0X1111000X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111100001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001000010000001  100000100X0011110");
    apply_vector ( 24'b001111100001000010000001,17'b100000100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001000010000001  0X1000100X1111111");
    apply_vector ( 24'b111111101001000010000001,17'b0X1000100X1111111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111100101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101000010000011  110100100X0111110");
    apply_vector ( 24'b010111100101000010000011,17'b110100100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101000010000001  0X1100100X0111110");
    apply_vector ( 24'b111111101101000010000001,17'b0X1100100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111100011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011000010000001  100010100X0111110");
    apply_vector ( 24'b001111100011000010000001,17'b100010100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011000010000001  0X1010100X0111110");
    apply_vector ( 24'b111111101011000010000001,17'b0X1010100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111100111000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111000010000000  110110100X0111110");
    apply_vector ( 24'b010111100111000010000000,17'b110110100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111101111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111000010000001  0X1110100X0111110");
    apply_vector ( 24'b111111101111000010000001,17'b0X1110100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000000010000001  101001000X0111110");
    apply_vector ( 24'b001100010000000010000001,17'b101001000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000000010000001  0X0101000X1XXXX01");
    apply_vector ( 24'b111100011000000010000001,17'b0X0101000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100000010000010  111101000X0XXXX00");
    apply_vector ( 24'b010100010100000010000010,17'b111101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100000010000000  0X0011000X0XXXX00");
    apply_vector ( 24'b111100011100000010000000,17'b0X0011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010000010000000  101011000X0XXXX00");
    apply_vector ( 24'b001100010010000010000000,17'b101011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010000010000000  0X0111000X0XXXX00");
    apply_vector ( 24'b111100011010000010000000,17'b0X0111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110000010000001  111111000X0XXXX00");
    apply_vector ( 24'b010100010110000010000001,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110000010000001  0X0000100X0XXXX00");
    apply_vector ( 24'b111100011110000010000001,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001000010000001  101000100X0XXXX00");
    apply_vector ( 24'b001100010001000010000001,17'b101000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001000010000001  0X0100100X1000111");
    apply_vector ( 24'b111100011001000010000001,17'b0X0100100X1000111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101000010000011  111100100X0000110");
    apply_vector ( 24'b010100010101000010000011,17'b111100100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101000010000000  0X0010100X0000110");
    apply_vector ( 24'b111100011101000010000000,17'b0X0010100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011000010000000  101010100X0000110");
    apply_vector ( 24'b001100010011000010000000,17'b101010100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011000010000000  0X0110100X0000110");
    apply_vector ( 24'b111100011011000010000000,17'b0X0110100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010100010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111000010000001  111110100X0000110");
    apply_vector ( 24'b010100010111000010000001,17'b111110100X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111000010000001  0X0001100X0000110");
    apply_vector ( 24'b111100011111000010000001,17'b0X0001100X0000110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000000010000001  100101000X0000110");
    apply_vector ( 24'b001110010000000010000001,17'b100101000X0000110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000000010000001  0X1101000X1XXXX01");
    apply_vector ( 24'b111110011000000010000001,17'b0X1101000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100000010000010  110011000X0XXXX00");
    apply_vector ( 24'b010110010100000010000010,17'b110011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100000010000001  0X1011000X0XXXX00");
    apply_vector ( 24'b111110011100000010000001,17'b0X1011000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110010010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010000010000000  100111000X0XXXX00");
    apply_vector ( 24'b001110010010000010000000,17'b100111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010000010000000  0X1111000X0XXXX00");
    apply_vector ( 24'b111110011010000010000000,17'b0X1111000X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110000010000001  110000100X0XXXX00");
    apply_vector ( 24'b010110010110000010000001,17'b110000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110000010000001  0X1000100X0XXXX00");
    apply_vector ( 24'b111110011110000010000001,17'b0X1000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001000010000001  100100100X0XXXX00");
    apply_vector ( 24'b001110010001000010000001,17'b100100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001000010000001  0X1100100X1XXXX01");
    apply_vector ( 24'b111110011001000010000001,17'b0X1100100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101000010000011  110010100X0XXXX00");
    apply_vector ( 24'b010110010101000010000011,17'b110010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101000010000001  0X1010100X0XXXX00");
    apply_vector ( 24'b111110011101000010000001,17'b0X1010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110010011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011000010000000  100110100X0XXXX00");
    apply_vector ( 24'b001110010011000010000000,17'b100110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011000010000000  0X1110100X0XXXX00");
    apply_vector ( 24'b111110011011000010000000,17'b0X1110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010110010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111000010000001  110001100X0XXXX00");
    apply_vector ( 24'b010110010111000010000001,17'b110001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111000010000001  0X1001100X0XXXX00");
    apply_vector ( 24'b111110011111000010000001,17'b0X1001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000000010000001  101101000X0XXXX00");
    apply_vector ( 24'b001101010000000010000001,17'b101101000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000000010000001  0X0011000X1101011");
    apply_vector ( 24'b111101011000000010000001,17'b0X0011000X1101011,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100000010000010  111011000X0101010");
    apply_vector ( 24'b010101010100000010000010,17'b111011000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100000010000000  0X0111000X0101010");
    apply_vector ( 24'b111101011100000010000000,17'b0X0111000X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010000010000001  101111000X0101010");
    apply_vector ( 24'b001101010010000010000001,17'b101111000X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010000010000000  0X0000100X0101010");
    apply_vector ( 24'b111101011010000010000000,17'b0X0000100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110000010000001  111000100X0101010");
    apply_vector ( 24'b010101010110000010000001,17'b111000100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110000010000001  0X0100100X0101010");
    apply_vector ( 24'b111101011110000010000001,17'b0X0100100X0101010,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001000010000001  101100100X0101010");
    apply_vector ( 24'b001101010001000010000001,17'b101100100X0101010,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001000010000001  0X0010100X1XXXX01");
    apply_vector ( 24'b111101011001000010000001,17'b0X0010100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101000010000011  111010100X0XXXX00");
    apply_vector ( 24'b010101010101000010000011,17'b111010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101011101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101000010000000  0X0110100X0XXXX00");
    apply_vector ( 24'b111101011101000010000000,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011000010000001  101110100X0XXXX00");
    apply_vector ( 24'b001101010011000010000001,17'b101110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011000010000000  0X0001100X0XXXX00");
    apply_vector ( 24'b111101011011000010000000,17'b0X0001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111000010000001  111001100X0XXXX00");
    apply_vector ( 24'b010101010111000010000001,17'b111001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111000010000001  0X0101100X0XXXX00");
    apply_vector ( 24'b111101011111000010000001,17'b0X0101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111010000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000000010000001  100011000X0XXXX00");
    apply_vector ( 24'b001111010000000010000001,17'b100011000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111011000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000000010000001  0X1011000X1011111");
    apply_vector ( 24'b111111011000000010000001,17'b0X1011000X1011111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111010100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100000010000010  110111000X0011110");
    apply_vector ( 24'b010111010100000010000010,17'b110111000X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100000010000001  0X1111000X0011110");
    apply_vector ( 24'b111111011100000010000001,17'b0X1111000X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111010010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010000010000001  100000100X0011110");
    apply_vector ( 24'b001111010010000010000001,17'b100000100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010000010000000  0X1000100X0011110");
    apply_vector ( 24'b111111011010000010000000,17'b0X1000100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111010110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110000010000001  110100100X0011110");
    apply_vector ( 24'b010111010110000010000001,17'b110100100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110000010000001  0X1100100X0011110");
    apply_vector ( 24'b111111011110000010000001,17'b0X1100100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111010001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001000010000001  100010100X0011110");
    apply_vector ( 24'b001111010001000010000001,17'b100010100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001000010000001  0X1010100X1101111");
    apply_vector ( 24'b111111011001000010000001,17'b0X1010100X1101111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111010101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101000010000011  110110100X0101110");
    apply_vector ( 24'b010111010101000010000011,17'b110110100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101000010000001  0X1110100X0101110");
    apply_vector ( 24'b111111011101000010000001,17'b0X1110100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111010011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011000010000001  100001100X0101110");
    apply_vector ( 24'b001111010011000010000001,17'b100001100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011000010000000  0X1001100X0101110");
    apply_vector ( 24'b111111011011000010000000,17'b0X1001100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111010111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111000010000001  110101100X0101110");
    apply_vector ( 24'b010111010111000010000001,17'b110101100X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111011111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111000010000001  0X1101100X0101110");
    apply_vector ( 24'b111111011111000010000001,17'b0X1101100X0101110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001100110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000000010000001  101011000X0101110");
    apply_vector ( 24'b001100110000000010000001,17'b101011000X0101110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111100111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000000010000001  0X0111000X1XXXX01");
    apply_vector ( 24'b111100111000000010000001,17'b0X0111000X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100000010000010  111111000X0XXXX00");
    apply_vector ( 24'b010100110100000010000010,17'b111111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100000010000000  0X0000100X0XXXX00");
    apply_vector ( 24'b111100111100000010000000,17'b0X0000100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010000010000000  101000100X0XXXX00");
    apply_vector ( 24'b001100110010000010000000,17'b101000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010000010000001  0X0100100X0XXXX00");
    apply_vector ( 24'b111100111010000010000001,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110000010000001  111100100X0XXXX00");
    apply_vector ( 24'b010100110110000010000001,17'b111100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110000010000001  0X0010100X0XXXX00");
    apply_vector ( 24'b111100111110000010000001,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001000010000001  101010100X0XXXX00");
    apply_vector ( 24'b001100110001000010000001,17'b101010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001000010000001  0X0110100X1XXXX01");
    apply_vector ( 24'b111100111001000010000001,17'b0X0110100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101000010000011  111110100X0XXXX00");
    apply_vector ( 24'b010100110101000010000011,17'b111110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101000010000000  0X0001100X0XXXX00");
    apply_vector ( 24'b111100111101000010000000,17'b0X0001100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001100110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011000010000000  101001100X0XXXX00");
    apply_vector ( 24'b001100110011000010000000,17'b101001100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011000010000001  0X0101100X0XXXX00");
    apply_vector ( 24'b111100111011000010000001,17'b0X0101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010100110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111000010000001  111101100X0XXXX00");
    apply_vector ( 24'b010100110111000010000001,17'b111101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111100111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111000010000001  0X0011100X0XXXX00");
    apply_vector ( 24'b111100111111000010000001,17'b0X0011100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001110110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000000010000001  100111000X0XXXX00");
    apply_vector ( 24'b001110110000000010000001,17'b100111000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111110111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000000010000001  0X1111000X1011111");
    apply_vector ( 24'b111110111000000010000001,17'b0X1111000X1011111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100000010000010  110000100X0011110");
    apply_vector ( 24'b010110110100000010000010,17'b110000100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100000010000001  0X1000100X0011110");
    apply_vector ( 24'b111110111100000010000001,17'b0X1000100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110110010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010000010000000  100100100X0011110");
    apply_vector ( 24'b001110110010000010000000,17'b100100100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010000010000001  0X1100100X0011110");
    apply_vector ( 24'b111110111010000010000001,17'b0X1100100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110000010000001  110010100X0011110");
    apply_vector ( 24'b010110110110000010000001,17'b110010100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110000010000001  0X1010100X0011110");
    apply_vector ( 24'b111110111110000010000001,17'b0X1010100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001000010000001  100110100X0011110");
    apply_vector ( 24'b001110110001000010000001,17'b100110100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001000010000001  0X1110100X1111111");
    apply_vector ( 24'b111110111001000010000001,17'b0X1110100X1111111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101000010000011  110001100X0111110");
    apply_vector ( 24'b010110110101000010000011,17'b110001100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101000010000001  0X1001100X0111110");
    apply_vector ( 24'b111110111101000010000001,17'b0X1001100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001110110011000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011000010000000  100101100X0111110");
    apply_vector ( 24'b001110110011000010000000,17'b100101100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011000010000001  0X1101100X0111110");
    apply_vector ( 24'b111110111011000010000001,17'b0X1101100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010110110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111000010000001  110011100X0111110");
    apply_vector ( 24'b010110110111000010000001,17'b110011100X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111110111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111000010000001  0X1011100X0111110");
    apply_vector ( 24'b111110111111000010000001,17'b0X1011100X0111110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000000010000001  101111000X0111110");
    apply_vector ( 24'b001101110000000010000001,17'b101111000X0111110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000000010000001  0X0000100X1XXXX01");
    apply_vector ( 24'b111101111000000010000001,17'b0X0000100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100000010000010  111000100X0XXXX00");
    apply_vector ( 24'b010101110100000010000010,17'b111000100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100000010000000  0X0100100X0XXXX00");
    apply_vector ( 24'b111101111100000010000000,17'b0X0100100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010000010000001  101100100X0XXXX00");
    apply_vector ( 24'b001101110010000010000001,17'b101100100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010000010000001  0X0010100X0XXXX00");
    apply_vector ( 24'b111101111010000010000001,17'b0X0010100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010101110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110000010000001  111010100X0XXXX00");
    apply_vector ( 24'b010101110110000010000001,17'b111010100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110000010000001  0X0110100X0XXXX00");
    apply_vector ( 24'b111101111110000010000001,17'b0X0110100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001101110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001000010000001  101110100X0XXXX00");
    apply_vector ( 24'b001101110001000010000001,17'b101110100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111101111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001000010000001  0X0001100X1011111");
    apply_vector ( 24'b111101111001000010000001,17'b0X0001100X1011111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101000010000011  111001100X0011110");
    apply_vector ( 24'b010101110101000010000011,17'b111001100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101000010000000  0X0101100X0011110");
    apply_vector ( 24'b111101111101000010000000,17'b0X0101100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001101110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011000010000001  101101100X0011110");
    apply_vector ( 24'b001101110011000010000001,17'b101101100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011000010000001  0X0011100X0011110");
    apply_vector ( 24'b111101111011000010000001,17'b0X0011100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010101110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111000010000001  111011100X0011110");
    apply_vector ( 24'b010101110111000010000001,17'b111011100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111101111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111000010000001  0X0111100X0011110");
    apply_vector ( 24'b111101111111000010000001,17'b0X0111100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111110000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000000010000001  100000100X0011110");
    apply_vector ( 24'b001111110000000010000001,17'b100000100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000000010000001  0X1000100X1011110");
    apply_vector ( 24'b111111111000000010000001,17'b0X1000100X1011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111110100000010000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100000010000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100000110000010  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100000110000010,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100000010000010  110100100X0011110");
    apply_vector ( 24'b010111110100000010000010,17'b110100100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111100000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100000010000001  0X1100100X0011110");
    apply_vector ( 24'b111111111100000010000001,17'b0X1100100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111110010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010000010000001  100010100X0011110");
    apply_vector ( 24'b001111110010000010000001,17'b100010100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111010000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010000010000001  0X1010100X0011110");
    apply_vector ( 24'b111111111010000010000001,17'b0X1010100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010111110110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110000010000001  110110100X0011110");
    apply_vector ( 24'b010111110110000010000001,17'b110110100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111110000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110000010000001  0X1110100X0011110");
    apply_vector ( 24'b111111111110000010000001,17'b0X1110100X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001111110001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001000010000001  100001100X0011110");
    apply_vector ( 24'b001111110001000010000001,17'b100001100X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111111111001000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001000010000001  0X1001100X1XXXX01");
    apply_vector ( 24'b111111111001000010000001,17'b0X1001100X1XXXX01,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111110101000010000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101000010000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101000110000011  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101000110000011,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101000010000011  110101100X0XXXX00");
    apply_vector ( 24'b010111110101000010000011,17'b110101100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111111101000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101000010000001  0X1101100X0XXXX00");
    apply_vector ( 24'b111111111101000010000001,17'b0X1101100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001111110011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011000010000001  100011100X0XXXX00");
    apply_vector ( 24'b001111110011000010000001,17'b100011100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111111011000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011000010000001  0X1011100X0XXXX00");
    apply_vector ( 24'b111111111011000010000001,17'b0X1011100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 010111110111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111000010000001  110111100X0XXXX00");
    apply_vector ( 24'b010111110111000010000001,17'b110111100X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111111111111000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111000010000001  0X1111100X0XXXX00");
    apply_vector ( 24'b111111111111000010000001,17'b0X1111100X0XXXX00,
                   24'b111111111111111111111111,17'b10111111101000011);
    $display ( "v 001000000000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000000010000001  100000000X0XXXX00");
    apply_vector ( 24'b001000000000000010000001,17'b100000000X0XXXX00,
                   24'b111111111111111111111111,17'b11111111101000011);
    $display ( "v 111000001000000010000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000000010000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000000110000001  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000000110000001,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000000010000001  0X1000000X1011111");
    apply_vector ( 24'b111000001000000010000001,17'b0X1000000X1011111,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000000100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100000010000000  110100000X0011110");
    apply_vector ( 24'b010000000100000010000000,17'b110100000X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000001100000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100000010000000  0X1100000X0011110");
    apply_vector ( 24'b111000001100000010000000,17'b0X1100000X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000000010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010000010000000  100010000X0011110");
    apply_vector ( 24'b001000000010000010000000,17'b100010000X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000001010000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010000010000000  0X1010000X0011110");
    apply_vector ( 24'b111000001010000010000000,17'b0X1010000X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000000110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110000010000000  110110000X0011110");
    apply_vector ( 24'b010000000110000010000000,17'b110110000X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000001110000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110000010000000  0X1110000X0011110");
    apply_vector ( 24'b111000001110000010000000,17'b0X1110000X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 001000000001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001000010000000  100001000X0011110");
    apply_vector ( 24'b001000000001000010000000,17'b100001000X0011110,
                   24'b111111111111111111111111,17'b11111111101111111);
    $display ( "v 111000001001000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001000010000000  0X1001000X0011110");
    apply_vector ( 24'b111000001001000010000000,17'b0X1001000X0011110,
                   24'b111111111111111111111111,17'b10111111101111111);
    $display ( "v 010000000101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101000110000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101000110000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101000010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000000101000010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001101000010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101000010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101100010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101100010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101000010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000001101000010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000000011011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000001011011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000000111011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000001111010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000010010000000  101000000X0XXXXX0");
    apply_vector ( 24'b001010000000010010000000,17'b101000000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000011010000000  0X0100000X0XXXXX0");
    apply_vector ( 24'b111010001000011010000000,17'b0X0100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100010010000000  111100000X0XXXXX0");
    apply_vector ( 24'b010010000100010010000000,17'b111100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100011010000000  0X0010010X0XXXXX0");
    apply_vector ( 24'b111010001100011010000000,17'b0X0010010X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010011010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001010000010011010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111010001010011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110011010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010010000110011010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111010001110011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001010010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010000001010010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010001001010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010000101011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010001101010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011011010000000  101011010X0XXXXX0");
    apply_vector ( 24'b001010000011011010000000,17'b101011010X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010001011011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010000111011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010001111011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000011010000000  100100000X0XXXXX0");
    apply_vector ( 24'b001001000000011010000000,17'b100100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000011010000000  0X1100000X0XXXXX0");
    apply_vector ( 24'b111001001000011010000000,17'b0X1100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100010010000000  110010000X0XXXXX0");
    apply_vector ( 24'b010001000100010010000000,17'b110010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100010010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111001001100010010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010011010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001001000010011010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010010010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111001001010010010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110011010000000  110001010X0XXXXX0");
    apply_vector ( 24'b010001000110011010000000,17'b110001010X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111001001110011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001000001011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001001001011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101011010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001000101011010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111001001101011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011011010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001000011011010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001001011010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001000111010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001001111011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000010010000000  101100000X0XXXXX0");
    apply_vector ( 24'b001011000000010010000000,17'b101100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000011010000000  0X0010010X0XXXXX0");
    apply_vector ( 24'b111011001000011010000000,17'b0X0010010X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100011010000000  111010000X0XXXXX0");
    apply_vector ( 24'b010011000100011010000000,17'b111010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111011001100011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010011010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001011000010011010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010010010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111011001010010010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110011010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010011000110011010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111011001110011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011000001011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011001001010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011000101010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111011001101011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011000011010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011011010000000  0X0000110X0XXXXX0");
    apply_vector ( 24'b111011001011011010000000,17'b0X0000110X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111011010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011000111011010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011001111011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000011010000000  100010000X0XXXXX0");
    apply_vector ( 24'b001000100000011010000000,17'b100010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000010010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111000101000010010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100010010000000  110110000X0XXXXX0");
    apply_vector ( 24'b010000100100010010000000,17'b110110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111000101100011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010011010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001000100010011010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111000101010011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110010010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000100110010010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000101110010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000100001011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000101001010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101011010000000  110111010X0XXXXX0");
    apply_vector ( 24'b010000100101011010000000,17'b110111010X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000101101011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001000100011011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111000101011011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111010010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010000100111010010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111000101111010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000011010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001010100000011010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111010101000011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100011010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010010100100011010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111010101100011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010010010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010100010010010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010101010010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010100110011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010101110010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001011010000000  101011010X0XXXXX0");
    apply_vector ( 24'b001010100001011010000000,17'b101011010X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010101001011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010100101011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010101101011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011010010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001010100011010010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111010101011010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111011010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010010100111011010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111010101111010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000011010000000  100110010X0XXXXX0");
    apply_vector ( 24'b001001100000011010000000,17'b100110010X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111001101000011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100011010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010001100100011010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100010010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111001101100010010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010010010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001100010010010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001101010011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110010010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001100110010010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110011010000000  0X1011010X0XXXXX0");
    apply_vector ( 24'b111001101110011010000000,17'b0X1011010X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001011010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001100001011010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001101001011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001100101011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001101101010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011010010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001001100011010010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111001101011011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111010010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010001100111010010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111011010000000  0X1010110X0XXXXX0");
    apply_vector ( 24'b111001101111011010000000,17'b0X1010110X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000011010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001011100000011010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111011101000011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100011010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010011100100011010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111011101100010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010010010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011100010010010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011101010011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011100110010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110011010000000  0X0111010X0XXXXX0");
    apply_vector ( 24'b111011101110011010000000,17'b0X0111010X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011100001010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011101001010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011100101010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011101101010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011010010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001011100011010010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111011101011010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111010010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010011100111010010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111011101111010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000010010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001000010000010010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000010010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111000011000010010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100010010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000010100010010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000011100010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000010010010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000011010010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110010010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000010110010010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000011110011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001010010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001000010001010010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111000011001010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101010010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010000010101010010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111000011101010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011010010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001000010011010010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111000011011010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111011010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010000010111011010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111000011111010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000010010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010010000010010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010011000010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100010010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010010100010010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010011100010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010010010010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010011010010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010010110011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010011110011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001010010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001010010001010010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111010011001010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101010010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010010010101010010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111010011101010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011010010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001010010011010010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111010011011011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111010010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010010010111010010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111010011111010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000010010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001010000010010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001011000010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100010010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001010100010010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111001011100010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001010010010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001011010011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001010110010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001011110011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001010010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001001010001010010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111001011001010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101010010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010001010101010010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111001011101010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011010010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001001010011010010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111001011011011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111011010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010001010111011010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111001011111010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000010010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011010000010010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011011000010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011010100010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111011011100010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011010010010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011011010011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110011010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011010110011010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011011110011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001010010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001011010001010010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111011011001010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101010010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010011010101010010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111011011101010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011011010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001011010011011010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111011011011010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111010010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010011010111010010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111011011111010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000110000010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000111000010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100010010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000110100010010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000111100010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001000110010011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111000111010010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110010010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010000110110010010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111000111110011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001010010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001000110001010010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111000111001010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101010010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010000110101010010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111000111101010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011011010000000  100001100X0XXXXX0");
    apply_vector ( 24'b001000110011011010000000,17'b100001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111000111011010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111011010000000  110101100X0XXXXX0");
    apply_vector ( 24'b010000110111011010000000,17'b110101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111010010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111000111111010010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010110000010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010111000010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010110100010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010111100010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001010110010011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111010111010010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110011010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010010110110011010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111010111110011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001010010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001010110001010010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111010111001010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101010010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010010110101010010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111010111101010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011011010000000  101001100X0XXXXX0");
    apply_vector ( 24'b001010110011011010000000,17'b101001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011011010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111010111011011010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111010010000000  111101100X0XXXXX0");
    apply_vector ( 24'b010010110111010010000000,17'b111101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111010010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111010111111010010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001110000010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001111000010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001110100010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001111100010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001001110010011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111001111010011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110010010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010001110110010010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111001111110011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001010010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001001110001010010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111001111001010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101010010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010001110101010010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111001111101010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011011010000000  100101100X0XXXXX0");
    apply_vector ( 24'b001001110011011010000000,17'b100101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011011010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111001111011011010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111011010000000  110011100X0XXXXX0");
    apply_vector ( 24'b010001110111011010000000,17'b110011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111010010000000  0X1011100X0XXXXX0");
    apply_vector ( 24'b111001111111010010000000,17'b0X1011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011110000010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011111000010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011110100010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011111100010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001011110010011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111011111010011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110011010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010011110110011010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111011111110011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001010010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001011110001010010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111011111001010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101010010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010011110101010010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101011010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111011111101011010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011010010000000  101101100X0XXXXX0");
    apply_vector ( 24'b001011110011010010000000,17'b101101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011010010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111011111011010010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111010010000000  111011100X0XXXXX0");
    apply_vector ( 24'b010011110111010010000000,17'b111011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111010010000000  0X0111100X0XXXXX0");
    apply_vector ( 24'b111011111111010010000000,17'b0X0111100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000010010000000  101000000X0XXXXX0");
    apply_vector ( 24'b001100000000010010000000,17'b101000000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000010010000000  0X0100000X0XXXXX0");
    apply_vector ( 24'b111100001000010010000000,17'b0X0100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100010010000000  111100000X0XXXXX0");
    apply_vector ( 24'b010100000100010010000000,17'b111100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100011010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111100001100011010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010010010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001100000010010010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010010010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111100001010010010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110010010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010100000110010010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111100001110011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001010010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001100000001010010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111100001001010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101010010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010100000101010010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111100001101011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100000011010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100001011010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100000111011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100001111010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000010010000000  100100000X0XXXXX0");
    apply_vector ( 24'b001110000000010010000000,17'b100100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000010010000000  0X1100000X0XXXXX0");
    apply_vector ( 24'b111110001000010010000000,17'b0X1100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100010010000000  110010000X0XXXXX0");
    apply_vector ( 24'b010110000100010010000000,17'b110010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100011010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111110001100011010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010010010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001110000010010010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010010010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111110001010010010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110011010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010110000110011010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111110001110011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001010010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001110000001010010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111110001001010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101010010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010110000101010010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111110001101011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110000011010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110001011011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110000111010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110001111010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000010010000000  101100000X0XXXXX0");
    apply_vector ( 24'b001101000000010010000000,17'b101100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000010010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111101001000010010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100010010000000  111010000X0XXXXX0");
    apply_vector ( 24'b010101000100010010000000,17'b111010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111101001100011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010010010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001101000010010010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111101001010011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110010010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010101000110010010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111101001110011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001010010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001101000001010010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111101001001010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010101000101010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111101001101011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101000011010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101001011011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111011010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101000111011010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101001111010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000010010000000  100010000X0XXXXX0");
    apply_vector ( 24'b001111000000010010000000,17'b100010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000010010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111111001000010010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100010010000000  110110000X0XXXXX0");
    apply_vector ( 24'b010111000100010010000000,17'b110110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111111001100011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010010010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001111000010010010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111111001010011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110011010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010111000110011010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111111001110011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001111000001010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111111001001010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101010010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010111000101010010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111111001101011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111000011011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111001011010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111010010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111000111010010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111001111010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000010010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001100100000010010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000010010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111100101000010010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100010010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010100100100010010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111100101100011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001100100010011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111100101010010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110010010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010100100110010010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111100101110011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100100001010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100101001010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100100101010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100101101011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001100100011011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111100101011010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111011010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010100100111011010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111100101111010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000010010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001110100000010010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000010010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111110101000010010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100010010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010110100100010010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111110101100011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001110100010011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111110101010010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110011010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010110100110011010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111110101110011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110100001010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110101001010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110100101010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110101101011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001110100011011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111110101011011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111010010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010110100111010010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111110101111010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000010010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001101100000010010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000010010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111101101000010010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100010010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010101100100010010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111101101100011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001101100010011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111101101010011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010101100110010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111101101110011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101100001010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101101001010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101100101010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101101101011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001101100011011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111101101011011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111011010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010101100111011010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111101101111010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000010010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001111100000010010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000010010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111111101000010010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100010010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010111100100010010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111111101100011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001111100010011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111111101010011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010111100110011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111111101110011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001010010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111100001010010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111101001010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111100101011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111101101010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011010010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001111100011010010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111111101011010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111010010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010111100111010010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111111101111010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000010010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001100010000010010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111100011000010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010100010100011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111100011100010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100010010010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100011010010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100010110010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100011110011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001010010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001100010001010010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111100011001010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101011010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010100010101011010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111100011101010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011010010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001100010011010010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111100011011010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111011010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010100010111011010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111100011111010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000010010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001110010000010010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111110011000010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100011010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010110010100011010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111110011100010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110010010010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110011010010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110010110011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110011110011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001010010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001110010001010010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111110011001010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101011010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010110010101011010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111110011101010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011010010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001110010011010010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111110011011011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111010010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010110010111010010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111110011111010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000010010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001101010000010010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111101011000010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100011010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010101010100011010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111101011100010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101010010010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101011010011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101010110010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101011110011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001010010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001101010001010010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111101011001010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101011010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010101010101011010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111101011101010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011010010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001101010011010010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011011010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111101011011011010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111011010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010101010111011010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111101011111010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001111010000010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111111011000010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010111010100011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111111011100010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010010010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111010010010010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111011010011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111010110011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111011110011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001010010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001111010001010010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111111011001010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101011010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010111010101011010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111111011101010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011011010000000  100001110X0XXXXX0");
    apply_vector ( 24'b001111010011011010000000,17'b100001110X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111111011011010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111010010000000  110101100X0XXXXX0");
    apply_vector ( 24'b010111010111010010000000,17'b110101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111010010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111111011111010010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100110000010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100111000010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100110100011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100111100010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001100110010011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111100111010010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110010010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010100110110010010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111100111110011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001010010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001100110001010010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111100111001010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101011010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010100110101011010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111100111101010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011011010000000  101001100X0XXXXX0");
    apply_vector ( 24'b001100110011011010000000,17'b101001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111100111011010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111011010000000  111101100X0XXXXX0");
    apply_vector ( 24'b010100110111011010000000,17'b111101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111010010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111100111111010010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110110000010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110111000010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110110100011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110111100010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001110110010011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111110111010010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110011010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010110110110011010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111110111110011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001010010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001110110001010010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111110111001010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101011010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010110110101011010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111110111101010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011011010000000  100101100X0XXXXX0");
    apply_vector ( 24'b001110110011011010000000,17'b100101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011011010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111110111011011010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111010010000000  110011100X0XXXXX0");
    apply_vector ( 24'b010110110111010010000000,17'b110011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111010010000000  0X1011100X0XXXXX0");
    apply_vector ( 24'b111110111111010010000000,17'b0X1011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101110000010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101111000010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100011010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101110100011010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101111100010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001101110010011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111101111010011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110010010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010101110110010010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111101111110011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001010010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001101110001010010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111101111001010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101011010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010101110101011010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111101111101010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011011010000000  101101100X0XXXXX0");
    apply_vector ( 24'b001101110011011010000000,17'b101101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011011010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111101111011011010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111011010000000  111011100X0XXXXX0");
    apply_vector ( 24'b010101110111011010000000,17'b111011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111010010000000  0X0111100X0XXXXX0");
    apply_vector ( 24'b111101111111010010000000,17'b0X0111100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000010010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111110000010010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111111000010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111110100011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111111100010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010011010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001111110010011010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111111111010011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110011010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010111110110011010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111111111110011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001010010000000  100001100X0XXXXX0");
    apply_vector ( 24'b001111110001010010000000,17'b100001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111111111001010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101011010000000  110101100X0XXXXX0");
    apply_vector ( 24'b010111110101011010000000,17'b110101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101011010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111111111101011010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011010010000000  100011100X0XXXXX0");
    apply_vector ( 24'b001111110011010010000000,17'b100011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011010010000000  0X1011100X0XXXXX0");
    apply_vector ( 24'b111111111011010010000000,17'b0X1011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111010010000000  110111100X0XXXXX0");
    apply_vector ( 24'b010111110111010010000000,17'b110111100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111010010000000  0X1111100X0XXXXX0");
    apply_vector ( 24'b111111111111010010000000,17'b0X1111100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000010010000000  100000000X0XXXXX0");
    apply_vector ( 24'b001000000000010010000000,17'b100000000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000010010000000  0X1000000X0XXXXX0");
    apply_vector ( 24'b111000001000010010000000,17'b0X1000000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100011010000000  110100000X0XXXXX0");
    apply_vector ( 24'b010000000100011010000000,17'b110100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100011010000000  0X1100000X0XXXXX0");
    apply_vector ( 24'b111000001100011010000000,17'b0X1100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010010010000000  100010000X0XXXXX0");
    apply_vector ( 24'b001000000010010010000000,17'b100010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010010010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111000001010010010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110010010000000  110110000X0XXXXX0");
    apply_vector ( 24'b010000000110010010000000,17'b110110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111000001110011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001010010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001000000001010010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001010010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111000001001010010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101011010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000000101011010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000001101011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000000011010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000001011010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000000111011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000001111010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000010010000000  101000000X0XXXXX0");
    apply_vector ( 24'b001010000000010010000000,17'b101000000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000010010000000  0X0100000X0XXXXX0");
    apply_vector ( 24'b111010001000010010000000,17'b0X0100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100011010000000  111100000X0XXXXX0");
    apply_vector ( 24'b010010000100011010000000,17'b111100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100011010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111010001100011010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010010010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001010000010010010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010010010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111010001010010010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110011010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010010000110011010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111010001110011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001010010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010000001010010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010001001010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010000101011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010001101011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010000011010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010001011011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010000111010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010001111010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000010010000000  100100000X0XXXXX0");
    apply_vector ( 24'b001001000000010010000000,17'b100100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000010010000000  0X1100000X0XXXXX0");
    apply_vector ( 24'b111001001000010010000000,17'b0X1100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100011010000000  110010000X0XXXXX0");
    apply_vector ( 24'b010001000100011010000000,17'b110010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100011010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111001001100011010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010010010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001001000010010010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111001001010011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110010010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010001000110010010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111001001110011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001010010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001000001010010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001001001010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101011010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001000101011010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111001001101011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001000011010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001001011011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001000111011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001001111010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000010010000000  101100000X0XXXXX0");
    apply_vector ( 24'b001011000000010010000000,17'b101100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000010010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111011001000010010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100011010000000  111010000X0XXXXX0");
    apply_vector ( 24'b010011000100011010000000,17'b111010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111011001100011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010010010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001011000010010010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111011001010011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110011010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010011000110011010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111011001110011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001010010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011000001010010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011001001010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101011010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011000101011010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111011001101011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011011010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011000011011010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011001011010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011000111010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011001111010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000010010000000  100010000X0XXXXX0");
    apply_vector ( 24'b001000100000010010000000,17'b100010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000010010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111000101000010010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100011010000000  110110000X0XXXXX0");
    apply_vector ( 24'b010000100100011010000000,17'b110110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111000101100011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010011010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001000100010011010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010010010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111000101010010010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110010010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000100110010010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000101110011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000100001010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000101001010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000100101011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000101101011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001000100011011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111000101011010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010000100111011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111000101111010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000010010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001010100000010010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000010010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111010101000010010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100011010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010010100100011010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111010101100011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010100010011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010101010010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010100110011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010101110011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010100001010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010101001010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010100101011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010101101011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001010100011011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111010101011011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111010010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010010100111010010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111010101111010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000010010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001001100000010010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000010010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111001101000010010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100011010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010001100100011010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111001101100011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001100010011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001101010011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110010010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001100110010010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111001101110011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001100001010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001101001010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001100101011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001101101011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001001100011011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111001101011011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111011010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010001100111011010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111001101111010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000010010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001011100000010010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000010010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111011101000010010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100011010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010011100100011010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111011101100011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011100010011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011101010011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110011010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011100110011010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111011101110011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011100001010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011101001011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011100101010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011101101010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011010010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001011100011010010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111011101011010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111010010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010011100111010010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111011101111010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000010010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001000010000010010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111000011000011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100010010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000010100010010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000011100010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000010010010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000011010010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110010010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000010110010010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000011110011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001010010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001000010001010010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111000011001011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101010010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010000010101010010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111000011101010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011010010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001000010011010010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111000011011010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111011010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010000010111011010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111000011111010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000010010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010010000010010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010011000011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100010010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010010100010010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010011100010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010010010010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010011010010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010010110011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010011110011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001010010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001010010001010010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111010011001011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101010010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010010010101010010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111010011101010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011010010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001010010011010010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111010011011011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111010010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010010010111010010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111010011111010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000010010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001010000010010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001011000011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100010010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001010100010010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111001011100010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001010010010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001011010011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001010110010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001011110011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001010010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001001010001010010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111001011001011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101010010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010001010101010010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111001011101010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011010010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001001010011010010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111001011011011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111011010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010001010111011010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111001011111010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000010010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011010000010010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011011000011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011010100010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111011011100010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011010010010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011011010011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110011010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011010110011010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011011110011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001010010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001011010001010010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111011011001011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101010010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010011010101010010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111011011101010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011011010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001011010011011010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111011011011010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111010010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010011010111010010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111011011111010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000110000010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000111000011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100010010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000110100010010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000111100010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001000110010011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111000111010010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110010010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010000110110010010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111000111110011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001010010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001000110001010010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111000111001011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101010010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010000110101010010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111000111101010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011011010000000  100001100X0XXXXX0");
    apply_vector ( 24'b001000110011011010000000,17'b100001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111000111011010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111011010000000  110101100X0XXXXX0");
    apply_vector ( 24'b010000110111011010000000,17'b110101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111010010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111000111111010010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010110000010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010111000011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010110100010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010111100010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001010110010011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111010111010010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110011010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010010110110011010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111010111110011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001010010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001010110001010010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111010111001011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101010010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010010110101010010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111010111101010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011011010000000  101001100X0XXXXX0");
    apply_vector ( 24'b001010110011011010000000,17'b101001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011011010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111010111011011010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111010010000000  111101100X0XXXXX0");
    apply_vector ( 24'b010010110111010010000000,17'b111101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111010010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111010111111010010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001110000010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001111000011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001110100010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001111100010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001001110010011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111001111010011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110010010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010001110110010010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111001111110011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001010010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001001110001010010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111001111001011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101010010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010001110101010010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111001111101010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011011010000000  100101100X0XXXXX0");
    apply_vector ( 24'b001001110011011010000000,17'b100101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011011010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111001111011011010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111011010000000  110011100X0XXXXX0");
    apply_vector ( 24'b010001110111011010000000,17'b110011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111010010000000  0X1011100X0XXXXX0");
    apply_vector ( 24'b111001111111010010000000,17'b0X1011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011110000010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011111000011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011110100010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011111100010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001011110010011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111011111010011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110011010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010011110110011010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111011111110011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001010010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001011110001010010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001011010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111011111001011010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101010010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010011110101010010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101011010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111011111101011010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011010010000000  101101100X0XXXXX0");
    apply_vector ( 24'b001011110011010010000000,17'b101101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011010010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111011111011010010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111010010000000  111011100X0XXXXX0");
    apply_vector ( 24'b010011110111010010000000,17'b111011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111010010000000  0X0111100X0XXXXX0");
    apply_vector ( 24'b111011111111010010000000,17'b0X0111100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000010010000000  101000000X0XXXXX0");
    apply_vector ( 24'b001100000000010010000000,17'b101000000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000011010000000  0X0100000X0XXXXX0");
    apply_vector ( 24'b111100001000011010000000,17'b0X0100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100010010000000  111100000X0XXXXX0");
    apply_vector ( 24'b010100000100010010000000,17'b111100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100011010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111100001100011010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010010010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001100000010010010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010010010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111100001010010010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110010010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010100000110010010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111100001110011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001010010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001100000001010010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111100001001011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101010010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010100000101010010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111100001101011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100000011010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100001011010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100000111011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100001111010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000010010000000  100100000X0XXXXX0");
    apply_vector ( 24'b001110000000010010000000,17'b100100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000011010000000  0X1100000X0XXXXX0");
    apply_vector ( 24'b111110001000011010000000,17'b0X1100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100010010000000  110010000X0XXXXX0");
    apply_vector ( 24'b010110000100010010000000,17'b110010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100011010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111110001100011010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010010010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001110000010010010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010010010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111110001010010010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110011010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010110000110011010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111110001110011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001010010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001110000001010010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111110001001011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101010010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010110000101010010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111110001101011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110000011010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110001011011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110000111010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110001111010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000010010000000  101100000X0XXXXX0");
    apply_vector ( 24'b001101000000010010000000,17'b101100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000011010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111101001000011010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100010010000000  111010000X0XXXXX0");
    apply_vector ( 24'b010101000100010010000000,17'b111010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111101001100011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010010010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001101000010010010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111101001010011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110010010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010101000110010010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111101001110011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001010010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001101000001010010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111101001001011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010101000101010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111101001101011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101000011010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101001011011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111011010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101000111011010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101001111010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000010010000000  100010000X0XXXXX0");
    apply_vector ( 24'b001111000000010010000000,17'b100010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000011010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111111001000011010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100010010000000  110110000X0XXXXX0");
    apply_vector ( 24'b010111000100010010000000,17'b110110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111111001100011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010010010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001111000010010010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111111001010011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110011010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010111000110011010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111111001110011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001111000001010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111111001001011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101010010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010111000101010010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111111001101011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111000011011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111001011010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111010010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111000111010010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111001111010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000010010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001100100000010010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111100101000011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100010010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010100100100010010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111100101100011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001100100010011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111100101010010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110010010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010100100110010010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111100101110011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100100001010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100101001011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100100101010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100101101011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001100100011011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111100101011010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111011010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010100100111011010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111100101111010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000010010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001110100000010010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111110101000011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100010010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010110100100010010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111110101100011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001110100010011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111110101010010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110011010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010110100110011010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111110101110011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110100001010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110101001011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110100101010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110101101011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001110100011011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111110101011011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111010010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010110100111010010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111110101111010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000010010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001101100000010010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111101101000011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100010010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010101100100010010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111101101100011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001101100010011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111101101010011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010101100110010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111101101110011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101100001010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101101001011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101100101010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101101101011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001101100011011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111101101011011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111011010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010101100111011010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111101101111010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000010010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001111100000010010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111111101000011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100010010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010111100100010010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100011010000000  0X1101010X0XXXXX0");
    apply_vector ( 24'b111111101100011010000000,17'b0X1101010X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001111100010011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111111101010011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010111100110011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111111101110011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001010010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111100001010010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111101001011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111100101011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111101101010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011010010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001111100011010010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111111101011010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111010010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010111100111010010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111111101111010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000010010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001100010000010010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111100011000011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010100010100011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111100011100010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100010010010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100011010010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100010110010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100011110011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001010010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001100010001010010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111100011001011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101011010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010100010101011010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111100011101010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011010010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001100010011010010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111100011011010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111011010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010100010111011010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111100011111010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000010010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001110010000010010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111110011000011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100011010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010110010100011010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111110011100010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110010010010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110011010010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110010110011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110011110011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001010010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001110010001010010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111110011001011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101011010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010110010101011010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111110011101010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011010010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001110010011010010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111110011011011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111010010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010110010111010010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111110011111010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000010010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001101010000010010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111101011000011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100011010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010101010100011010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111101011100010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101010010010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101011010011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101010110010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101011110011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001010010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001101010001010010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111101011001011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101011010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010101010101011010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111101011101010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011010010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001101010011010010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011011010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111101011011011010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111011010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010101010111011010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111101011111010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001111010000010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111111011000011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010111010100011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111111011100010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010010010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111010010010010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111011010011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111010110011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111011110011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001010010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001111010001010010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111111011001011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101011010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010111010101011010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111111011101010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011011010000000  100001100X0XXXXX0");
    apply_vector ( 24'b001111010011011010000000,17'b100001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111111011011010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111010010000000  110101100X0XXXXX0");
    apply_vector ( 24'b010111010111010010000000,17'b110101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111010010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111111011111010010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100110000010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100111000011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100110100011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100111100010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001100110010011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111100111010010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110010010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010100110110010010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111100111110011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001010010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001100110001010010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111100111001011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101011010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010100110101011010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111100111101010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011011010000000  101001100X0XXXXX0");
    apply_vector ( 24'b001100110011011010000000,17'b101001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111100111011010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111011010000000  111101100X0XXXXX0");
    apply_vector ( 24'b010100110111011010000000,17'b111101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111010010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111100111111010010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110110000010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110111000011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110110100011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110111100010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001110110010011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111110111010010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110011010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010110110110011010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111110111110011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001010010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001110110001010010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111110111001011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101011010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010110110101011010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111110111101010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011011010000000  100101100X0XXXXX0");
    apply_vector ( 24'b001110110011011010000000,17'b100101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011011010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111110111011011010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111010010000000  110011100X0XXXXX0");
    apply_vector ( 24'b010110110111010010000000,17'b110011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111010010000000  0X1011100X0XXXXX0");
    apply_vector ( 24'b111110111111010010000000,17'b0X1011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101110000010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101111000011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100011010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101110100011010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101111100010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001101110010011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111101111010011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110010010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010101110110010010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111101111110011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001010010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001101110001010010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001011010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111101111001011010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101011010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010101110101011010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111101111101010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011011010000000  101101100X0XXXXX0");
    apply_vector ( 24'b001101110011011010000000,17'b101101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011011010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111101111011011010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111011010000000  111011100X0XXXXX0");
    apply_vector ( 24'b010101110111011010000000,17'b111011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111010010000000  0X0111100X0XXXXX0");
    apply_vector ( 24'b111101111111010010000000,17'b0X0111100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000010010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111110000010010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111111000011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111110100011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111111100010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010011010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001111110010011010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111111111010011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110011010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010111110110011010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111111111110011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001010010000000  100001100X0XXXXX0");
    apply_vector ( 24'b001111110001010010000000,17'b100001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001011010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111111111001011010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101011010000000  110101100X0XXXXX0");
    apply_vector ( 24'b010111110101011010000000,17'b110101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101011010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111111111101011010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011010010000000  100011100X0XXXXX0");
    apply_vector ( 24'b001111110011010010000000,17'b100011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011010010000000  0X1011100X0XXXXX0");
    apply_vector ( 24'b111111111011010010000000,17'b0X1011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111010010000000  110111100X0XXXXX0");
    apply_vector ( 24'b010111110111010010000000,17'b110111100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111010010000000  0X1111100X0XXXXX0");
    apply_vector ( 24'b111111111111010010000000,17'b0X1111100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000010010000000  100000000X0XXXXX0");
    apply_vector ( 24'b001000000000010010000000,17'b100000000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000011010000000  0X1000000X0XXXXX0");
    apply_vector ( 24'b111000001000011010000000,17'b0X1000000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100011010000000  110100000X0XXXXX0");
    apply_vector ( 24'b010000000100011010000000,17'b110100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100011010000000  0X1100000X0XXXXX0");
    apply_vector ( 24'b111000001100011010000000,17'b0X1100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010010010000000  100010000X0XXXXX0");
    apply_vector ( 24'b001000000010010010000000,17'b100010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010010010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111000001010010010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110010010000000  110110000X0XXXXX0");
    apply_vector ( 24'b010000000110010010000000,17'b110110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111000001110011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001010010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001000000001010010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111000001001011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101011010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000000101011010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000001101011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000000011010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000001011010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000000111011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000001111010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000010010000000  101000000X0XXXXX0");
    apply_vector ( 24'b001010000000010010000000,17'b101000000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000011010000000  0X0100000X0XXXXX0");
    apply_vector ( 24'b111010001000011010000000,17'b0X0100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100011010000000  111100000X0XXXXX0");
    apply_vector ( 24'b010010000100011010000000,17'b111100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100011010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111010001100011010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010010010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001010000010010010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010010010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111010001010010010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110011010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010010000110011010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111010001110011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001010010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010000001010010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010001001011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010000101011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010001101011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010000011010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010001011011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010000111010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010001111010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000010010000000  100100000X0XXXXX0");
    apply_vector ( 24'b001001000000010010000000,17'b100100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000011010000000  0X1100000X0XXXXX0");
    apply_vector ( 24'b111001001000011010000000,17'b0X1100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100011010000000  110010000X0XXXXX0");
    apply_vector ( 24'b010001000100011010000000,17'b110010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100011010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111001001100011010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010010010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001001000010010010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111001001010011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110010010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010001000110010010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111001001110011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001010010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001000001010010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001001001011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101011010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001000101011010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111001001101011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001000011010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001001011011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001000111011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001001111010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000010010000000  101100000X0XXXXX0");
    apply_vector ( 24'b001011000000010010000000,17'b101100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000011010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111011001000011010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100011010000000  111010000X0XXXXX0");
    apply_vector ( 24'b010011000100011010000000,17'b111010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111011001100011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010010010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001011000010010010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111011001010011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110011010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010011000110011010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111011001110011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001010010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011000001010010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011001001011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101011010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011000101011010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111011001101011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011011010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011000011011010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011001011010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011000111010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011001111010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000010010000000  100010000X0XXXXX0");
    apply_vector ( 24'b001000100000010010000000,17'b100010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000011010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111000101000011010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100011010000000  110110000X0XXXXX0");
    apply_vector ( 24'b010000100100011010000000,17'b110110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111000101100011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010011010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001000100010011010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010010010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111000101010010010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110010010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000100110010010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000101110011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000100001010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001011010000000  0X1011010X0XXXXX0");
    apply_vector ( 24'b111000101001011010000000,17'b0X1011010X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000100101011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000101101011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001000100011011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111000101011010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010000100111011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111000101111010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000010010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001010100000010010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111010101000011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100011010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010010100100011010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111010101100011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010100010011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010101010010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010100110011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010101110011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010100001010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010101001011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010100101011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010101101011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001010100011011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111010101011011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111010010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010010100111010010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111010101111010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000010010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001001100000010010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111001101000011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100011010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010001100100011010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111001101100011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001100010011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001101010011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110010010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001100110010010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111001101110011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001100001010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001101001011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001100101011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001101101011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001001100011011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111001101011011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111011010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010001100111011010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111001101111010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000010010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001011100000010010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111011101000011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100011010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010011100100011010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111011101100011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011100010011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011101010011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110011010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011100110011010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111011101110011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001011010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011100001011010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011101001010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011100101010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011101101010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011010010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001011100011010010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111011101011010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111010010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010011100111010010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111011101111010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000011010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001000010000011010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000010010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111000011000010010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100010010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000010100010010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000011100010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000010010010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000011010010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110010010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000010110010010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000011110011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001000010001011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111000011001010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101010010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010000010101010010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111000011101010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011010010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001000010011010010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111000011011010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111011010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010000010111011010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111000011111010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010010000011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010011000010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100010010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010010100010010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010011100010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010010010010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010011010010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010010110011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010011110011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001010010001011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111010011001010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101010010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010010010101010010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111010011101010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011010010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001010010011010010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111010011011011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111010010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010010010111010010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111010011111010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001010000011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001011000010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100010010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001010100010010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111001011100010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001010010010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001011010011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001010110010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001011110011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001001010001011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111001011001010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101010010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010001010101010010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111001011101010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011010010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001001010011010010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111001011011011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111011010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010001010111011010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111001011111010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011010000011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011011000010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011010100010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111011011100010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011010010010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011011010011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110011010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011010110011010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011011110011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001011010001011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111011011001010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101010010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010011010101010010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111011011101010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011011010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001011010011011010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111011011011010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111010010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010011010111010010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111011011111010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000110000011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000111000010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100010010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000110100010010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000111100010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001000110010011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111000111010010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110010010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010000110110010010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111000111110011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001011010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001000110001011010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111000111001010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101010010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010000110101010010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111000111101010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011011010000000  100001100X0XXXXX0");
    apply_vector ( 24'b001000110011011010000000,17'b100001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111000111011010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111011010000000  110101100X0XXXXX0");
    apply_vector ( 24'b010000110111011010000000,17'b110101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111010010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111000111111010010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000011010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010110000011010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010111000010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010110100010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010111100010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001010110010011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111010111010010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110011010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010010110110011010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111010111110011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001011010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001010110001011010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111010111001010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101010010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010010110101010010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111010111101010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011011010000000  101001100X0XXXXX0");
    apply_vector ( 24'b001010110011011010000000,17'b101001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011011010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111010111011011010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111010010000000  111101100X0XXXXX0");
    apply_vector ( 24'b010010110111010010000000,17'b111101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111010010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111010111111010010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000011010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001110000011010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001111000010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001110100010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001111100010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001001110010011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111001111010011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110010010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010001110110010010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111001111110011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001011010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001001110001011010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111001111001010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101010010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010001110101010010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111001111101010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011011010000000  100101100X0XXXXX0");
    apply_vector ( 24'b001001110011011010000000,17'b100101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011011010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111001111011011010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111011010000000  110011100X0XXXXX0");
    apply_vector ( 24'b010001110111011010000000,17'b110011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111010010000000  0X1011100X0XXXXX0");
    apply_vector ( 24'b111001111111010010000000,17'b0X1011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000011010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011110000011010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011111000010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011110100010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011111100010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001011110010011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111011111010011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110011010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010011110110011010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111011111110011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001011010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001011110001011010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111011111001010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101010010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010011110101010010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101011010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111011111101011010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011010010000000  101101100X0XXXXX0");
    apply_vector ( 24'b001011110011010010000000,17'b101101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011010010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111011111011010010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111010010000000  111011100X0XXXXX0");
    apply_vector ( 24'b010011110111010010000000,17'b111011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111010010000000  0X0111100X0XXXXX0");
    apply_vector ( 24'b111011111111010010000000,17'b0X0111100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000011010000000  101000000X0XXXXX0");
    apply_vector ( 24'b001100000000011010000000,17'b101000000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000010010000000  0X0100000X0XXXXX0");
    apply_vector ( 24'b111100001000010010000000,17'b0X0100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100010010000000  111100000X0XXXXX0");
    apply_vector ( 24'b010100000100010010000000,17'b111100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100011010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111100001100011010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010010010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001100000010010010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010010010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111100001010010010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110010010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010100000110010010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111100001110011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001100000001011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111100001001010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101010010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010100000101010010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111100001101011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100000011010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100001011010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100000111011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100001111010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000011010000000  100100000X0XXXXX0");
    apply_vector ( 24'b001110000000011010000000,17'b100100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000010010000000  0X1100000X0XXXXX0");
    apply_vector ( 24'b111110001000010010000000,17'b0X1100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100010010000000  110010000X0XXXXX0");
    apply_vector ( 24'b010110000100010010000000,17'b110010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100011010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111110001100011010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010010010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001110000010010010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010010010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111110001010010010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110011010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010110000110011010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111110001110011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001110000001011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111110001001010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101010010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010110000101010010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111110001101011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110000011010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011011010000000  0X1111010X0XXXXX0");
    apply_vector ( 24'b111110001011011010000000,17'b0X1111010X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110000111010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110001111010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000011010000000  101100000X0XXXXX0");
    apply_vector ( 24'b001101000000011010000000,17'b101100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000010010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111101001000010010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100010010000000  111010000X0XXXXX0");
    apply_vector ( 24'b010101000100010010000000,17'b111010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111101001100011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010010010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001101000010010010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111101001010011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110010010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010101000110010010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111101001110011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001101000001011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111101001001010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010101000101010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111101001101011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101000011010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101001011011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111011010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101000111011010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101001111010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000011010000000  100010000X0XXXXX0");
    apply_vector ( 24'b001111000000011010000000,17'b100010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000010010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111111001000010010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100010010000000  110110000X0XXXXX0");
    apply_vector ( 24'b010111000100010010000000,17'b110110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111111001100011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010010010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001111000010010010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111111001010011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110011010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010111000110011010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111111001110011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001111000001011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111111001001010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101010010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010111000101010010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111111001101011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111000011011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111001011010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111010010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111000111010010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111001111010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000011010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001100100000011010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000010010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111100101000010010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100010010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010100100100010010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111100101100011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001100100010011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111100101010010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110010010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010100100110010010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111100101110011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001011010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100100001011010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100101001010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100100101010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100101101011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001100100011011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111100101011010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111011010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010100100111011010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111100101111010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000011010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001110100000011010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000010010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111110101000010010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100010010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010110100100010010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111110101100011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001110100010011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111110101010010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110011010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010110100110011010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111110101110011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001011010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110100001011010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110101001010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110100101010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110101101011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001110100011011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111110101011011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111010010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010110100111010010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111110101111010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000011010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001101100000011010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000010010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111101101000010010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100010010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010101100100010010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111101101100011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001101100010011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111101101010011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010101100110010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111101101110011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001011010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101100001011010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101101001010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101100101010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101101101011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001101100011011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111101101011011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111011010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010101100111011010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111101101111010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000011010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001111100000011010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000010010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111111101000010010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100010010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010111100100010010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111111101100011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001111100010011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111111101010011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010111100110011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111111101110011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111100001011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111101001010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111100101011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111101101010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011010010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001111100011010010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111111101011010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111010010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010111100111010010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111111101111010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001100010000011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111100011000010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010100010100011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111100011100010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100010010010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100011010010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100010110010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100011110011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001100010001011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111100011001010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101011010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010100010101011010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111100011101010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011010010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001100010011010010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111100011011010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111011010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010100010111011010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111100011111010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001110010000011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111110011000010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100011010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010110010100011010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111110011100010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110010010010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110011010010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110010110011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110011110011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001110010001011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111110011001010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101011010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010110010101011010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111110011101010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011010010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001110010011010010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111110011011011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111010010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010110010111010010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111110011111010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001101010000011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111101011000010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100011010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010101010100011010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111101011100010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101010010010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101011010011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101010110010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101011110011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001101010001011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111101011001010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101011010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010101010101011010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111101011101010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011010010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001101010011010010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011011010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111101011011011010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111011010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010101010111011010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111101011111010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001111010000011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111111011000010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010111010100011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111111011100010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010010010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111010010010010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111011010011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111010110011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111011110011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001011010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001111010001011010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111111011001010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101011010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010111010101011010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111111011101010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011011010000000  100001100X0XXXXX0");
    apply_vector ( 24'b001111010011011010000000,17'b100001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111111011011010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111010010000000  110101100X0XXXXX0");
    apply_vector ( 24'b010111010111010010000000,17'b110101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111010010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111111011111010010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000011010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100110000011010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100111000010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100110100011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100111100010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001100110010011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111100111010010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110010010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010100110110010010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111100111110011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001011010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001100110001011010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111100111001010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101011010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010100110101011010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111100111101010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011011010000000  101001100X0XXXXX0");
    apply_vector ( 24'b001100110011011010000000,17'b101001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111100111011010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111011010000000  111101100X0XXXXX0");
    apply_vector ( 24'b010100110111011010000000,17'b111101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111010010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111100111111010010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000011010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110110000011010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110111000010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110110100011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110111100010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001110110010011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111110111010010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110011010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010110110110011010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111110111110011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001011010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001110110001011010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111110111001010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101011010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010110110101011010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111110111101010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011011010000000  100101100X0XXXXX0");
    apply_vector ( 24'b001110110011011010000000,17'b100101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011011010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111110111011011010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111010010000000  110011100X0XXXXX0");
    apply_vector ( 24'b010110110111010010000000,17'b110011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111010010000000  0X1011100X0XXXXX0");
    apply_vector ( 24'b111110111111010010000000,17'b0X1011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000011010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101110000011010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101111000010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100011010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101110100011010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101111100010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001101110010011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111101111010011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110010010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010101110110010010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111101111110011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001011010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001101110001011010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111101111001010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101011010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010101110101011010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111101111101010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011011010000000  101101100X0XXXXX0");
    apply_vector ( 24'b001101110011011010000000,17'b101101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011011010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111101111011011010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111011010000000  111011100X0XXXXX0");
    apply_vector ( 24'b010101110111011010000000,17'b111011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111010010000000  0X0111100X0XXXXX0");
    apply_vector ( 24'b111101111111010010000000,17'b0X0111100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111110000011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111111000010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111110100011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111111100010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010011010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001111110010011010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111111111010011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110011010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010111110110011010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111111111110011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001011010000000  100001100X0XXXXX0");
    apply_vector ( 24'b001111110001011010000000,17'b100001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111111111001010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101011010000000  110101100X0XXXXX0");
    apply_vector ( 24'b010111110101011010000000,17'b110101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101011010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111111111101011010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011010010000000  100011100X0XXXXX0");
    apply_vector ( 24'b001111110011010010000000,17'b100011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011010010000000  0X1011100X0XXXXX0");
    apply_vector ( 24'b111111111011010010000000,17'b0X1011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111010010000000  110111100X0XXXXX0");
    apply_vector ( 24'b010111110111010010000000,17'b110111100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111010010000000  0X1111100X0XXXXX0");
    apply_vector ( 24'b111111111111010010000000,17'b0X1111100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000011010000000  100000000X0XXXXX0");
    apply_vector ( 24'b001000000000011010000000,17'b100000000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000010010000000  0X1000000X0XXXXX0");
    apply_vector ( 24'b111000001000010010000000,17'b0X1000000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100011010000000  110100000X0XXXXX0");
    apply_vector ( 24'b010000000100011010000000,17'b110100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100011010000000  0X1100000X0XXXXX0");
    apply_vector ( 24'b111000001100011010000000,17'b0X1100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010010010000000  100010000X0XXXXX0");
    apply_vector ( 24'b001000000010010010000000,17'b100010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010010010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111000001010010010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110010010000000  110110000X0XXXXX0");
    apply_vector ( 24'b010000000110010010000000,17'b110110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111000001110011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001011010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001000000001011010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001010010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111000001001010010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101011010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000000101011010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000001101011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000000011010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000001011010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000000111011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000001111010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000011010000000  101000000X0XXXXX0");
    apply_vector ( 24'b001010000000011010000000,17'b101000000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000010010000000  0X0100000X0XXXXX0");
    apply_vector ( 24'b111010001000010010000000,17'b0X0100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100011010000000  111100000X0XXXXX0");
    apply_vector ( 24'b010010000100011010000000,17'b111100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100011010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111010001100011010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010010010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001010000010010010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010010010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111010001010010010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110011010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010010000110011010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111010001110011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010000001011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010001001010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010000101011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010001101011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010000011010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010001011011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010000111010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010001111010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000011010000000  100100000X0XXXXX0");
    apply_vector ( 24'b001001000000011010000000,17'b100100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000010010000000  0X1100000X0XXXXX0");
    apply_vector ( 24'b111001001000010010000000,17'b0X1100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100011010000000  110010000X0XXXXX0");
    apply_vector ( 24'b010001000100011010000000,17'b110010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100011010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111001001100011010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010010010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001001000010010010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111001001010011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110010010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010001000110010010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111001001110011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001000001011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001001001010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101011010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001000101011010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111001001101011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001000011010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001001011011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001000111011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001001111010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000011010000000  101100000X0XXXXX0");
    apply_vector ( 24'b001011000000011010000000,17'b101100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000010010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111011001000010010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100011010000000  111010000X0XXXXX0");
    apply_vector ( 24'b010011000100011010000000,17'b111010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111011001100011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010010010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001011000010010010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111011001010011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110011010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010011000110011010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111011001110011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011000001011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011001001010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101011010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011000101011010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111011001101011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011011010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011000011011010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011001011010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011000111010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011001111010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000011010000000  100010000X0XXXXX0");
    apply_vector ( 24'b001000100000011010000000,17'b100010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000010010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111000101000010010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100011010000000  110110000X0XXXXX0");
    apply_vector ( 24'b010000100100011010000000,17'b110110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111000101100011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010011010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001000100010011010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010010010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111000101010010010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110010010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000100110010010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000101110011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000100001011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000101001010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000100101011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000101101011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001000100011011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111000101011010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010000100111011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111000101111010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000011010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001010100000011010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000010010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111010101000010010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100011010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010010100100011010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111010101100011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010100010011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010101010010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010100110011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010101110011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001011010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010100001011010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010101001010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010100101011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010101101011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001010100011011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111010101011011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111010010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010010100111010010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111010101111010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000011010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001001100000011010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000010010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111001101000010010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100011010000000  110001010X0XXXXX0");
    apply_vector ( 24'b010001100100011010000000,17'b110001010X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111001101100011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001100010011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001101010011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110010010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001100110010010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111001101110011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001011010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001100001011010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101001010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001101001010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001100101011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001101101011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001001100011011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111001101011011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111011010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010001100111011010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111001101111010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000011010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001011100000011010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101000010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000010010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111011101000010010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100011010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010011100100011010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111011101100011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011100010011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011101010011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110011010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011100110011010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111011101110011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100001011010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011100001011010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101001011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011101001011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100101010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011100101010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101101010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011101101010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100011010010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001011100011010010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101011010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111011101011010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100111010010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010011100111010010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101111010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111011101111010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010000011010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001000010000011010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011000011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111000011000011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010100010010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000010100010010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011100010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000011100010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010010010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000010010010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011010010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000011010010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010110010010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000010110010010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011110011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000011110011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010001011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001000010001011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011001011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111000011001011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010101010010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010000010101010010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011101010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111000011101010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000010011010010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001000010011010010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011011010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111000011011010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000010111011010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010000010111011010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000011111010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111000011111010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010000011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010010000011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011000011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010011000011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010100010010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010010100010010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011100010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010011100010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010010010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010010010010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011010010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010011010010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010110011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010010110011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011110011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010011110011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010001011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001010010001011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011001011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111010011001011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010101010010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010010010101010010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011101010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111010011101010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010010011010010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001010010011010010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011011011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111010011011011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010010111010010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010010010111010010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010011111010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111010011111010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010000011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001010000011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011000011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001011000011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010100010010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001010100010010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011100010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111001011100010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010010010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001010010010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011010011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001011010011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010110010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001010110010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011110011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001011110011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010001011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001001010001011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011001011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111001011001011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010101010010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010001010101010010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011101010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111001011101010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001010011010010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001001010011010010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011011011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111001011011011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001010111011010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010001010111011010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001011111010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111001011111010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010000011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011010000011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011000011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011011000011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010100010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011010100010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011100010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111011011100010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010010010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011010010010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011010011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011011010011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010110011010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011010110011010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011110011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011011110011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010001011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001011010001011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011001011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111011011001011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010101010010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010011010101010010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011101010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111011011101010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011010011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011010011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011010011011010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001011010011011010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011011010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111011011011010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011010111010010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010011010111010010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011011111010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111011011111010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110000011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000110000011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111000011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000111000011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110100010010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000110100010010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111100010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000111100010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110010011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001000110010011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111010010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111000111010010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110110010010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010000110110010010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111110011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111000111110011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110001011010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001000110001011010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111001011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111000111001011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110101010010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010000110101010010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111101010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111000111101010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000110011011010000000  100001100X0XXXXX0");
    apply_vector ( 24'b001000110011011010000000,17'b100001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111011010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111000111011010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000110111011010000000  110101110X0XXXXX0");
    apply_vector ( 24'b010000110111011010000000,17'b110101110X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000111111010010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111000111111010010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110000011010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010110000011010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111000011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010111000011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110100010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010110100010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111100010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010111100010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110010011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001010110010011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111010010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111010111010010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110110011010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010010110110011010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111110011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111010111110011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110001011010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001010110001011010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111001011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111010111001011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110101010010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010010110101010010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111101010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111010111101010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010110011011010000000  101001100X0XXXXX0");
    apply_vector ( 24'b001010110011011010000000,17'b101001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111011011010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111010111011011010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010110111010010000000  111101100X0XXXXX0");
    apply_vector ( 24'b010010110111010010000000,17'b111101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010111111010010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111010111111010010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110000011010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001110000011010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111000011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001111000011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110100010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001110100010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111100010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001111100010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110010011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001001110010011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111010011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111001111010011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110110010010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010001110110010010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111110011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111001111110011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110001011010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001001110001011010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111001011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111001111001011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110101010010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010001110101010010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111101010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111001111101010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001110011011010000000  100101100X0XXXXX0");
    apply_vector ( 24'b001001110011011010000000,17'b100101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111011011010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111001111011011010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001110111011010000000  110011100X0XXXXX0");
    apply_vector ( 24'b010001110111011010000000,17'b110011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001111111010010000000  0X1011100X0XXXXX0");
    apply_vector ( 24'b111001111111010010000000,17'b0X1011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110000011010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011110000011010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111000011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011111000011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110100010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011110100010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111100010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011111100010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110010011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001011110010011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111010011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111011111010011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110110011010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010011110110011010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111110011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111011111110011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110001011010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001011110001011010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111001011010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111011111001011010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110101010010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010011110101010010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111101011010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111011111101011010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011110011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011110011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011110011010010000000  101101100X0XXXXX0");
    apply_vector ( 24'b001011110011010010000000,17'b101101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111011010010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111011111011010010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011110111010010000000  111011100X0XXXXX0");
    apply_vector ( 24'b010011110111010010000000,17'b111011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011111111010010000000  0X0111100X0XXXXX0");
    apply_vector ( 24'b111011111111010010000000,17'b0X0111100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000000011010000000  101000000X0XXXXX0");
    apply_vector ( 24'b001100000000011010000000,17'b101000000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001000011010000000  0X0100000X0XXXXX0");
    apply_vector ( 24'b111100001000011010000000,17'b0X0100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000100010010000000  111100000X0XXXXX0");
    apply_vector ( 24'b010100000100010010000000,17'b111100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001100011010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111100001100011010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000010010010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001100000010010010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001010010010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111100001010010010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000110010010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010100000110010010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001110011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111100001110011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000001011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001100000001011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001001011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111100001001011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000101010010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010100000101010010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001101011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111100001101011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100000011010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100000011010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001011010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100001011010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100000111011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100000111011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100001111010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100001111010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000000011010000000  100100000X0XXXXX0");
    apply_vector ( 24'b001110000000011010000000,17'b100100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001000011010000000  0X1100000X0XXXXX0");
    apply_vector ( 24'b111110001000011010000000,17'b0X1100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000100010010000000  110010000X0XXXXX0");
    apply_vector ( 24'b010110000100010010000000,17'b110010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001100011010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111110001100011010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000010010010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001110000010010010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001010010010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111110001010010010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000110011010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010110000110011010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001110011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111110001110011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000001011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001110000001011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001001011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111110001001011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000101010010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010110000101010010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001101011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111110001101011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110000011010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110000011010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001011011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110001011011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110000111010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110000111010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110001111010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110001111010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000000011010000000  101100000X0XXXXX0");
    apply_vector ( 24'b001101000000011010000000,17'b101100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001000011010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111101001000011010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000100010010000000  111010000X0XXXXX0");
    apply_vector ( 24'b010101000100010010000000,17'b111010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001100011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111101001100011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000010010010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001101000010010010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001010011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111101001010011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000110010010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010101000110010010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001110011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111101001110011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000001011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001101000001011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001001011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111101001001011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000101010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010101000101010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001101011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111101001101011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101000011010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101000011010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001011011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101001011011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101000111011010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101000111011010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101001111010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101001111010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000000011010000000  100010000X0XXXXX0");
    apply_vector ( 24'b001111000000011010000000,17'b100010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001000011010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111111001000011010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000100010010000000  110110000X0XXXXX0");
    apply_vector ( 24'b010111000100010010000000,17'b110110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001100011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111111001100011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000010010010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001111000010010010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001010011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111111001010011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000110011010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010111000110011010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001110011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111111001110011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000001011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001111000001011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001001011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111111001001011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000101010010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010111000101010010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001101011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111111001101011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111000011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111000011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111000011011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111000011011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001011010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111001011010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111000111010010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111000111010010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111001111010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111001111010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100000011010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001100100000011010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101000011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111100101000011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100100010010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010100100100010010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101100011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111100101100011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100010011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001100100010011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101010010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111100101010010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100110010010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010100100110010010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101110011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111100101110011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100001011010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100100001011010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101001011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100101001011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100101010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100100101010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101101011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100101101011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100100011011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001100100011011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101011010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111100101011010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100100111011010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010100100111011010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100101111010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111100101111010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100000011010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001110100000011010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101000011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111110101000011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100100010010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010110100100010010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101100011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111110101100011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100010011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001110100010011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101010010010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111110101010010010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100110011010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010110100110011010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101110011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111110101110011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100001011010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110100001011010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101001011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110101001011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100101010010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110100101010010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101101011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110101101011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110100011011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001110100011011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101011011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111110101011011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110100111010010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010110100111010010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110101111010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111110101111010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100000011010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001101100000011010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101000011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111101101000011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100100010010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010101100100010010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101100011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111101101100011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100010011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001101100010011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101010011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111101101010011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100110010010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010101100110010010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101110011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111101101110011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100001011010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101100001011010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101001011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101101001011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100101010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101100101010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101101011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101101101011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101100011011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001101100011011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101011011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111101101011011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101100111011010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010101100111011010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101101111010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111101101111010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100000011010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001111100000011010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101000011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111111101000011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100100010010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010111100100010010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101100011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111111101100011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100010011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001111100010011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101010011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111111101010011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100110011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010111100110011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101110011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111111101110011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100001011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111100001011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101001011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111101001011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100101011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111100101011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101101010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111101101010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111100011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111100011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111100011010010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001111100011010010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101011010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111111101011010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111100111010010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010111100111010010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111101111010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111111101111010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010000011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001100010000011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011000011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111100011000011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010100011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010100010100011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011100010010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111100011100010010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010010010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100010010010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011010010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100011010010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010110010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100010110010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011110011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100011110011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010001011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001100010001011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011001011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111100011001011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010101011010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010100010101011010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011101010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111100011101010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100010011010010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001100010011010010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011011010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111100011011010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100010111011010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010100010111011010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100011111010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111100011111010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010000011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001110010000011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011000011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111110011000011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010100011010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010110010100011010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011100010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111110011100010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010010010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110010010010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011010010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110011010010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010110011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110010110011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011110011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110011110011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010001011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001110010001011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011001011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111110011001011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010101011010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010110010101011010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011101010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111110011101010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110010011010010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001110010011010010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011011011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111110011011011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110010111010010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010110010111010010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110011111010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111110011111010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010000011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001101010000011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011000011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111101011000011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010100011010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010101010100011010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011100010010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111101011100010010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010010010010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101010010010010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011010011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101011010011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010110010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101010110010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011110011010000000  0X0100110X0XXXXX0");
    apply_vector ( 24'b111101011110011010000000,17'b0X0100110X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010001011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001101010001011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011001011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111101011001011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010101011010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010101010101011010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011101010010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111101011101010010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101010011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101010011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101010011010010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001101010011010010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011011011010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111101011011011010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101010111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101010111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101010111011010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010101010111011010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101011111010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111101011111010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010000011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001111010000011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011000011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111111011000011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010100011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010111010100011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011100010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111111011100010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010010010010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111010010010010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011010011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111011010011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010110011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111010110011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011110011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111011110011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010001011010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001111010001011010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011001011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111111011001011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010101011010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010111010101011010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011101010010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111111011101010010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111010011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111010011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111010011011010000000  100001100X0XXXXX0");
    apply_vector ( 24'b001111010011011010000000,17'b100001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011011010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111111011011010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111010111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111010111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111010111010010000000  110101100X0XXXXX0");
    apply_vector ( 24'b010111010111010010000000,17'b110101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111011111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111011111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111011111010010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111111011111010010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110000011010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001100110000011010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111000011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111100111000011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110100011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010100110100011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111100010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111100111100010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110010011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001100110010011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111010010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111100111010010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110110010010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010100110110010010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111110011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111100111110011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110001011010000000  101010100X0XXXXX0");
    apply_vector ( 24'b001100110001011010000000,17'b101010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111001011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111100111001011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110101011010000000  111110100X0XXXXX0");
    apply_vector ( 24'b010100110101011010000000,17'b111110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111101010010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111100111101010010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001100110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001100110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001100110011011010000000  101001100X0XXXXX0");
    apply_vector ( 24'b001100110011011010000000,17'b101001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111011010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111100111011010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010100110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010100110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010100110111011010000000  111101100X0XXXXX0");
    apply_vector ( 24'b010100110111011010000000,17'b111101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111100111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111100111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111100111111010010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111100111111010010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110000011010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001110110000011010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111000011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111110111000011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110100011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010110110100011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111100010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111110111100010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110010011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001110110010011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111010010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111110111010010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110110011010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010110110110011010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111110011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111110111110011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110001011010000000  100110100X0XXXXX0");
    apply_vector ( 24'b001110110001011010000000,17'b100110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111001011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111110111001011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110101011010000000  110001100X0XXXXX0");
    apply_vector ( 24'b010110110101011010000000,17'b110001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111101010010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111110111101010010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001110110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001110110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001110110011011010000000  100101100X0XXXXX0");
    apply_vector ( 24'b001110110011011010000000,17'b100101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111011011010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111110111011011010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010110110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010110110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010110110111010010000000  110011100X0XXXXX0");
    apply_vector ( 24'b010110110111010010000000,17'b110011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111110111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111110111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111110111111010010000000  0X1011100X0XXXXX0");
    apply_vector ( 24'b111110111111010010000000,17'b0X1011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110000011010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001101110000011010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111000011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111101111000011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110100011010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010101110100011010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111100010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111101111100010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110010011010000000  101100100X0XXXXX0");
    apply_vector ( 24'b001101110010011010000000,17'b101100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111010011010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111101111010011010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110110010010000000  111010100X0XXXXX0");
    apply_vector ( 24'b010101110110010010000000,17'b111010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111110011010000000  0X0110100X0XXXXX0");
    apply_vector ( 24'b111101111110011010000000,17'b0X0110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110001011010000000  101110100X0XXXXX0");
    apply_vector ( 24'b001101110001011010000000,17'b101110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111001011010000000  0X0001100X0XXXXX0");
    apply_vector ( 24'b111101111001011010000000,17'b0X0001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110101011010000000  111001100X0XXXXX0");
    apply_vector ( 24'b010101110101011010000000,17'b111001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111101010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111101110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111101010010000000  0X0101100X0XXXXX0");
    apply_vector ( 24'b111101111101010010000000,17'b0X0101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001101110011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001101110011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001101110011011010000000  101101100X0XXXXX0");
    apply_vector ( 24'b001101110011011010000000,17'b101101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111011011010000000  0X0011100X0XXXXX0");
    apply_vector ( 24'b111101111011011010000000,17'b0X0011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010101110111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010101110111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010101110111011010000000  111011100X0XXXXX0");
    apply_vector ( 24'b010101110111011010000000,17'b111011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111101111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111101111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111101111111010010000000  0X0111100X0XXXXX0");
    apply_vector ( 24'b111101111111010010000000,17'b0X0111100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110000011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001111110000011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111000011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111111111000011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110100011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010111110100011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111100010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111100110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111100010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111111111100010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110010011010000000  100010100X0XXXXX0");
    apply_vector ( 24'b001111110010011010000000,17'b100010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111010011010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111111111010011010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110110011010000000  110110100X0XXXXX0");
    apply_vector ( 24'b010111110110011010000000,17'b110110100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111110011010000000  0X1110100X0XXXXX0");
    apply_vector ( 24'b111111111110011010000000,17'b0X1110100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110001011010000000  100001100X0XXXXX0");
    apply_vector ( 24'b001111110001011010000000,17'b100001100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111001011010000000  0X1001100X0XXXXX0");
    apply_vector ( 24'b111111111001011010000000,17'b0X1001100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110101011010000000  110101100X0XXXXX0");
    apply_vector ( 24'b010111110101011010000000,17'b110101100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111101011010000000  0X1101100X0XXXXX0");
    apply_vector ( 24'b111111111101011010000000,17'b0X1101100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001111110011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001111110011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001111110011010010000000  100011100X0XXXXX0");
    apply_vector ( 24'b001111110011010010000000,17'b100011100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111011010010000000  0X1011100X0XXXXX0");
    apply_vector ( 24'b111111111011010010000000,17'b0X1011100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010111110111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010111110111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010111110111010010000000  110111100X0XXXXX0");
    apply_vector ( 24'b010111110111010010000000,17'b110111100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111111111111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111111111111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111111111111010010000000  0X1111100X0XXXXX0");
    apply_vector ( 24'b111111111111010010000000,17'b0X1111100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000000011010000000  100000000X0XXXXX0");
    apply_vector ( 24'b001000000000011010000000,17'b100000000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001000011010000000  0X1000000X0XXXXX0");
    apply_vector ( 24'b111000001000011010000000,17'b0X1000000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000100011010000000  110100000X0XXXXX0");
    apply_vector ( 24'b010000000100011010000000,17'b110100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001100011010000000  0X1100000X0XXXXX0");
    apply_vector ( 24'b111000001100011010000000,17'b0X1100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000010010010000000  100010000X0XXXXX0");
    apply_vector ( 24'b001000000010010010000000,17'b100010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001010010010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111000001010010010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000110010010000000  110110000X0XXXXX0");
    apply_vector ( 24'b010000000110010010000000,17'b110110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001110011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111000001110011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000001011010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001000000001011010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001001011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111000001001011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000101011010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000000101011010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001101011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000001101011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000000011010010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000000011010010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001011010010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000001011010010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000000111011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000000111011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000001111010010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000001111010010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000000011010000000  101000010X0XXXXX0");
    apply_vector ( 24'b001010000000011010000000,17'b101000010X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001000011010000000  0X0100000X0XXXXX0");
    apply_vector ( 24'b111010001000011010000000,17'b0X0100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000100011010000000  111100000X0XXXXX0");
    apply_vector ( 24'b010010000100011010000000,17'b111100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001100011010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111010001100011010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000010010010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001010000010010010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001010010010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111010001010010010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000110011010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010010000110011010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001110011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111010001110011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000001011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010000001011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001001011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010001001011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000101011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010000101011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001101011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010001101011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010000011010010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010000011010010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001011011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010001011011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010000111010010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010000111010010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010001111010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010001111010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000000011010000000  100100000X0XXXXX0");
    apply_vector ( 24'b001001000000011010000000,17'b100100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001000011010000000  0X1100000X0XXXXX0");
    apply_vector ( 24'b111001001000011010000000,17'b0X1100000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000100011010000000  110010000X0XXXXX0");
    apply_vector ( 24'b010001000100011010000000,17'b110010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001100011010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111001001100011010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000010010010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001001000010010010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001010011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111001001010011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000110010010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010001000110010010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001110011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111001001110011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000001011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001000001011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001001011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001001001011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000101011010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001000101011010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001101011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111001001101011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001000011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001000011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001000011010010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001000011010010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001011011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001001011011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001000111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001000111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001000111011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001000111011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001001111010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001001111010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000000011010000000  101100000X0XXXXX0");
    apply_vector ( 24'b001011000000011010000000,17'b101100000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001000011010000000  0X0010000X0XXXXX0");
    apply_vector ( 24'b111011001000011010000000,17'b0X0010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000100011010000000  111010000X0XXXXX0");
    apply_vector ( 24'b010011000100011010000000,17'b111010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001100011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111011001100011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000010010010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001011000010010010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001010011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111011001010011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000110011010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010011000110011010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001110011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111011001110011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000001011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011000001011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001001011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011001001011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000101011010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011000101011010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001101011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111011001101011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011000011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011000011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011000011011010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011000011011010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001011010010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011001011010010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011000111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011000111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011000111010010000000  111000100X0XXXXX0");
    apply_vector ( 24'b010011000111010010000000,17'b111000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011001111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011001111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011001111010010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111011001111010010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100000011010000000  100010000X0XXXXX0");
    apply_vector ( 24'b001000100000011010000000,17'b100010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101000011010000000  0X1010000X0XXXXX0");
    apply_vector ( 24'b111000101000011010000000,17'b0X1010000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100100011010000000  110110000X0XXXXX0");
    apply_vector ( 24'b010000100100011010000000,17'b110110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101100011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111000101100011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100010011010000000  100001000X0XXXXX0");
    apply_vector ( 24'b001000100010011010000000,17'b100001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101010010010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111000101010010010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100110010010000000  110101000X0XXXXX0");
    apply_vector ( 24'b010000100110010010000000,17'b110101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101110011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111000101110011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100001011010000000  100011000X0XXXXX0");
    apply_vector ( 24'b001000100001011010000000,17'b100011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101001011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111000101001011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100101011010000000  110111000X0XXXXX0");
    apply_vector ( 24'b010000100101011010000000,17'b110111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101101011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111000101101011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001000100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001000100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001000100011011010000000  100000100X0XXXXX0");
    apply_vector ( 24'b001000100011011010000000,17'b100000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101011010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101011110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101011010010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111000101011010010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010000100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010000100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010000100111011010000000  110100100X0XXXXX0");
    apply_vector ( 24'b010000100111011010000000,17'b110100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111000101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111000101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111000101111010010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111000101111010010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100000011010000000  101010000X0XXXXX0");
    apply_vector ( 24'b001010100000011010000000,17'b101010000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101000011010000000  0X0110000X0XXXXX0");
    apply_vector ( 24'b111010101000011010000000,17'b0X0110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100100011010000000  111110000X0XXXXX0");
    apply_vector ( 24'b010010100100011010000000,17'b111110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101100011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111010101100011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100010011010000000  101001000X0XXXXX0");
    apply_vector ( 24'b001010100010011010000000,17'b101001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101010010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101010110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101010010010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111010101010010010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100110011010000000  111101000X0XXXXX0");
    apply_vector ( 24'b010010100110011010000000,17'b111101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101110011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111010101110011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100001011010000000  101011000X0XXXXX0");
    apply_vector ( 24'b001010100001011010000000,17'b101011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101001011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111010101001011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100101011010000000  111111000X0XXXXX0");
    apply_vector ( 24'b010010100101011010000000,17'b111111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101101011010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111010101101011010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001010100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001010100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001010100011011010000000  101000100X0XXXXX0");
    apply_vector ( 24'b001010100011011010000000,17'b101000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101011011010000000  0X0100100X0XXXXX0");
    apply_vector ( 24'b111010101011011010000000,17'b0X0100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010010100111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010010100111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010010100111010010000000  111100100X0XXXXX0");
    apply_vector ( 24'b010010100111010010000000,17'b111100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111010101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111010101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111010101111010010000000  0X0010100X0XXXXX0");
    apply_vector ( 24'b111010101111010010000000,17'b0X0010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100000011010000000  100110000X0XXXXX0");
    apply_vector ( 24'b001001100000011010000000,17'b100110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101000011010000000  0X1110000X0XXXXX0");
    apply_vector ( 24'b111001101000011010000000,17'b0X1110000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100100011010000000  110001000X0XXXXX0");
    apply_vector ( 24'b010001100100011010000000,17'b110001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101100011010000000  0X1001000X0XXXXX0");
    apply_vector ( 24'b111001101100011010000000,17'b0X1001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100010011010000000  100101000X0XXXXX0");
    apply_vector ( 24'b001001100010011010000000,17'b100101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101010011010000000  0X1101000X0XXXXX0");
    apply_vector ( 24'b111001101010011010000000,17'b0X1101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100110010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100110110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100110010010000000  110011000X0XXXXX0");
    apply_vector ( 24'b010001100110010010000000,17'b110011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101110011010000000  0X1011000X0XXXXX0");
    apply_vector ( 24'b111001101110011010000000,17'b0X1011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100001011010000000  100111000X0XXXXX0");
    apply_vector ( 24'b001001100001011010000000,17'b100111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101001011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101001111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101001011010000000  0X1111000X0XXXXX0");
    apply_vector ( 24'b111001101001011010000000,17'b0X1111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100101011010000000  110000100X0XXXXX0");
    apply_vector ( 24'b010001100101011010000000,17'b110000100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101101011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101101111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101101011010000000  0X1000100X0XXXXX0");
    apply_vector ( 24'b111001101101011010000000,17'b0X1000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001001100011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001001100011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001001100011011010000000  100100100X0XXXXX0");
    apply_vector ( 24'b001001100011011010000000,17'b100100100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101011011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101011111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101011011010000000  0X1100100X0XXXXX0");
    apply_vector ( 24'b111001101011011010000000,17'b0X1100100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010001100111011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010001100111111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010001100111011010000000  110010100X0XXXXX0");
    apply_vector ( 24'b010001100111011010000000,17'b110010100X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111001101111010010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111010010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111110010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111001101111110010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111001101111010010000000  0X1010100X0XXXXX0");
    apply_vector ( 24'b111001101111010010000000,17'b0X1010100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100000011010000000  101110000X0XXXXX0");
    apply_vector ( 24'b001011100000011010000000,17'b101110000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101000011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101000111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101000011010000000  0X0001000X0XXXXX0");
    apply_vector ( 24'b111011101000011010000000,17'b0X0001000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100100011010000000  111001000X0XXXXX0");
    apply_vector ( 24'b010011100100011010000000,17'b111001000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101100011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101100111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101100011010000000  0X0101000X0XXXXX0");
    apply_vector ( 24'b111011101100011010000000,17'b0X0101000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b001011100010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 001011100010011010000000  101101000X0XXXXX0");
    apply_vector ( 24'b001011100010011010000000,17'b101101000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101010011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101010111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101010011010000000  0X0011000X0XXXXX0");
    apply_vector ( 24'b111011101010011010000000,17'b0X0011000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 010011100110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b010011100110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 010011100110011010000000  111011000X0XXXXX0");
    apply_vector ( 24'b010011100110011010000000,17'b111011000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101110011010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110011010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110111010000000  XXXXXXXXXXXXXXXXX");
    apply_vector ( 24'b111011101110111010000000,17'bXXXXXXXXXXXXXXXXX,
                   24'b111111111111111111111111,17'b00000000000000000);
    $display ( "v 111011101110011010000000  0X0111000X0XXXXX0");
    apply_vector ( 24'b111011101110011010000000,17'b0X0111000X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    $display ( "v 001011100001000010000000  101111000X0XXXXX0");
    apply_vector ( 24'b001011100001000010000000,17'b101111000X0XXXXX0,
                   24'b111111111111111111111111,17'b11111111101000001);
    $display ( "v 111011101001000010000000  0X0000100X0XXXXX0");
    apply_vector ( 24'b111011101001000010000000,17'b0X0000100X0XXXXX0,
                   24'b111111111111111111111111,17'b10111111101000001);
    if ( errors == 0 )
      begin
        $display( "Simulation OK" );
        $display( "All vectors passed" );
      end
    else
      begin
        $display( "" );
        $display( "Simulation Failed" );
        $display( "" );
        if (  errors_Q0 > 0 )
          $display ( "       ", errors_Q0, " errors with Q0",) ;
        if (  errors_Q1 > 0 )
          $display ( "       ", errors_Q1, " errors with Q1",) ;
        if (  errors_Q3 > 0 )
          $display ( "       ", errors_Q3, " errors with Q3",) ;
        if (  errors_Q4 > 0 )
          $display ( "       ", errors_Q4, " errors with Q4",) ;
        if (  errors_Q5 > 0 )
          $display ( "       ", errors_Q5, " errors with Q5",) ;
        if (  errors_Q6 > 0 )
          $display ( "       ", errors_Q6, " errors with Q6",) ;
        if (  errors_Q7 > 0 )
          $display ( "       ", errors_Q7, " errors with Q7",) ;
        if (  errors_Q12 > 0 )
          $display ( "       ", errors_Q12, " errors with Q12",) ;
        if (  errors_Q15 > 0 )
          $display ( "       ", errors_Q15, " errors with Q15",) ;
        if (  errors_Q16 > 0 )
          $display ( "       ", errors_Q16, " errors with Q16",) ;
        if (  errors_Q17 > 0 )
          $display ( "       ", errors_Q17, " errors with Q17",) ;
        if (  errors_Q18 > 0 )
          $display ( "       ", errors_Q18, " errors with Q18",) ;
        if (  errors_Q19 > 0 )
          $display ( "       ", errors_Q19, " errors with Q19",) ;
        if (  errors_Q20 > 0 )
          $display ( "       ", errors_Q20, " errors with Q20",) ;
        if (  errors_Q21 > 0 )
          $display ( "       ", errors_Q21, " errors with Q21",) ;
        if (  errors_Q22 > 0 )
          $display ( "       ", errors_Q22, " errors with Q22",) ;
        if (  errors_Q23 > 0 )
          $display ( "       ", errors_Q23, " errors with Q23",) ;
        $display( "" );
        $display( "Total: ", errors, " errors");
        $display( "" );
      end
    $stop;
    $finish;
  end

// function declaration

task apply_vector;

  input [23:0] stimulus_vector;
  input [16:0] expected_vector;
  input [23:0] stimulus_mask;
  input [16:0] expected_mask;

  begin
    `ifdef set_x_to_0
      {A0,A1,A2,A3,A4,A5,A6,A7,A8,A9,A10,A11,A12,A13,A14,A15,A16,A17,A18,A19,A20,A21,A22,A23} = stimulus_vector & stimulus_mask ;
    `else
      {A0,A1,A2,A3,A4,A5,A6,A7,A8,A9,A10,A11,A12,A13,A14,A15,A16,A17,A18,A19,A20,A21,A22,A23} = stimulus_vector;
    `endif
    #500
    check_vector( expected_vector, expected_mask );
    #500
    $display("");
  end

endtask
task check_vector;

  input [16:0] expected_vector;
  input [16:0] mask_vector;

  reg [16:0] received_vector;
  reg [16:0] difference_vector;

  integer local_errors;

  begin
    local_errors = 0;
    received_vector = {Q0,Q1,Q3,Q4,Q5,Q6,Q7,Q12,Q15,Q16,Q17,Q18,Q19,Q20,Q21,Q22,Q23};
    difference_vector = ( received_vector ^ expected_vector ) & mask_vector ;
    $display( "r                           %b", received_vector );
    $display( "                            %s", error_point( difference_vector ) );
    if ( expected_vector[16] !== 1'bX )
      if ( expected_vector[16] !== Q0)
        begin
          $display( "error with Q0 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q0 = errors_Q0 + 1;
        end
    if ( expected_vector[15] !== 1'bX )
      if ( expected_vector[15] !== Q1)
        begin
          $display( "error with Q1 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q1 = errors_Q1 + 1;
        end
    if ( expected_vector[14] !== 1'bX )
      if ( expected_vector[14] !== Q3)
        begin
          $display( "error with Q3 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q3 = errors_Q3 + 1;
        end
    if ( expected_vector[13] !== 1'bX )
      if ( expected_vector[13] !== Q4)
        begin
          $display( "error with Q4 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q4 = errors_Q4 + 1;
        end
    if ( expected_vector[12] !== 1'bX )
      if ( expected_vector[12] !== Q5)
        begin
          $display( "error with Q5 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q5 = errors_Q5 + 1;
        end
    if ( expected_vector[11] !== 1'bX )
      if ( expected_vector[11] !== Q6)
        begin
          $display( "error with Q6 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q6 = errors_Q6 + 1;
        end
    if ( expected_vector[10] !== 1'bX )
      if ( expected_vector[10] !== Q7)
        begin
          $display( "error with Q7 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q7 = errors_Q7 + 1;
        end
    if ( expected_vector[9] !== 1'bX )
      if ( expected_vector[9] !== Q12)
        begin
          $display( "error with Q12 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q12 = errors_Q12 + 1;
        end
    if ( expected_vector[8] !== 1'bX )
      if ( expected_vector[8] !== Q15)
        begin
          $display( "error with Q15 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q15 = errors_Q15 + 1;
        end
    if ( expected_vector[7] !== 1'bX )
      if ( expected_vector[7] !== Q16)
        begin
          $display( "error with Q16 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q16 = errors_Q16 + 1;
        end
    if ( expected_vector[6] !== 1'bX )
      if ( expected_vector[6] !== Q17)
        begin
          $display( "error with Q17 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q17 = errors_Q17 + 1;
        end
    if ( expected_vector[5] !== 1'bX )
      if ( expected_vector[5] !== Q18)
        begin
          $display( "error with Q18 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q18 = errors_Q18 + 1;
        end
    if ( expected_vector[4] !== 1'bX )
      if ( expected_vector[4] !== Q19)
        begin
          $display( "error with Q19 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q19 = errors_Q19 + 1;
        end
    if ( expected_vector[3] !== 1'bX )
      if ( expected_vector[3] !== Q20)
        begin
          $display( "error with Q20 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q20 = errors_Q20 + 1;
        end
    if ( expected_vector[2] !== 1'bX )
      if ( expected_vector[2] !== Q21)
        begin
          $display( "error with Q21 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q21 = errors_Q21 + 1;
        end
    if ( expected_vector[1] !== 1'bX )
      if ( expected_vector[1] !== Q22)
        begin
          $display( "error with Q22 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q22 = errors_Q22 + 1;
        end
    if ( expected_vector[0] !== 1'bX )
      if ( expected_vector[0] !== Q23)
        begin
          $display( "error with Q23 @ %d ns", $time );
          local_errors = local_errors + 1;
          errors_Q23 = errors_Q23 + 1;
        end
    if ( local_errors > 0 ) $display( "" );
    errors = errors + local_errors;
  end

endtask
function [135:0] error_point;

  input [16:0] in_vector;
  integer i, j;
  begin
    error_point[ 7 : 0 ] = ( in_vector[ 0 ] === 0 ) ? " " : "^";
    error_point[ 15 : 8 ] = ( in_vector[ 1 ] === 0 ) ? " " : "^";
    error_point[ 23 : 16 ] = ( in_vector[ 2 ] === 0 ) ? " " : "^";
    error_point[ 31 : 24 ] = ( in_vector[ 3 ] === 0 ) ? " " : "^";
    error_point[ 39 : 32 ] = ( in_vector[ 4 ] === 0 ) ? " " : "^";
    error_point[ 47 : 40 ] = ( in_vector[ 5 ] === 0 ) ? " " : "^";
    error_point[ 55 : 48 ] = ( in_vector[ 6 ] === 0 ) ? " " : "^";
    error_point[ 63 : 56 ] = ( in_vector[ 7 ] === 0 ) ? " " : "^";
    error_point[ 71 : 64 ] = ( in_vector[ 8 ] === 0 ) ? " " : "^";
    error_point[ 79 : 72 ] = ( in_vector[ 9 ] === 0 ) ? " " : "^";
    error_point[ 87 : 80 ] = ( in_vector[ 10 ] === 0 ) ? " " : "^";
    error_point[ 95 : 88 ] = ( in_vector[ 11 ] === 0 ) ? " " : "^";
    error_point[ 103 : 96 ] = ( in_vector[ 12 ] === 0 ) ? " " : "^";
    error_point[ 111 : 104 ] = ( in_vector[ 13 ] === 0 ) ? " " : "^";
    error_point[ 119 : 112 ] = ( in_vector[ 14 ] === 0 ) ? " " : "^";
    error_point[ 127 : 120 ] = ( in_vector[ 15 ] === 0 ) ? " " : "^";
    error_point[ 135 : 128 ] = ( in_vector[ 16 ] === 0 ) ? " " : "^";
  end

endfunction


endmodule

